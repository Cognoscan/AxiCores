/**
# PS7 Wrapper #

Wraps the PS7 primitive using SystemVerilog Interfaces, making for a much more 
manageable netlist.

Although the port list is more compact, it is still recommended that a shim 
module be used, such that the rest of the system only sees the necessary ports. 
An example is included as ps7_shim.sv.
*/

///////////////////////////////////////////////////////////////////////////
// Module Declaration {{{
///////////////////////////////////////////////////////////////////////////
module ps7_wrapper
(
    // Dedicated PS Signal Pins
    inout logic PS_CLK,
    inout logic PS_POR_B,
    inout logic PS_SRST_B,
    ddr_if.controller ddr,
    inout  wire [53:0] MIO,

    // FCLK
    output logic [3:0] fclk_CLK,      ///< Generated clocks for use by FPGA logic
    input  logic [3:0] fclk_CLKTRIGN, ///< Disables related clock if set (may not be implemented)
    output logic [3:0] fclk_RESETN,   ///< Asynchronous resets loosely related to FCLK outputs

    /// Central Interconnect Clock Disable
    input  logic FPGAIDLEN, ///< Assert to let central interconnect clocks to shut off is all conditions are met

    // EVENT
    output logic [1:0] event_STANDBYWFE, ///< Asserted when CPU waiting for an event
    output logic [1:0] event_STANDBYWFI, ///< Asserted when CPU waiting for interrupt
    input  logic event_EVENTI,           ///< Causes CPUs to wake from WFE state
    output logic event_EVENTO,           ///< Asserted when a CPU has exectued the SEV instruction

    // AXI3 Bus Masters
    axi3_if.master m_axi_gp0, ///< Master GP0 - 32-bit data, 32-bit address, 12-bit ID
    axi3_if.master m_axi_gp1, ///< Master GP0 - 32-bit data, 32-bit address, 12-bit ID

    // AXI3 ACP Bus Slave
    axi3_if.slave s_axi_acp,             ///< Slave ACP - 64-bit data, 32-bit address, 3-bit ID
    input  logic [4:0] s_axi_acp_awuser, ///< Slave ACP - User pins to inform Snoop Control Unit
    input  logic [4:0] s_axi_acp_aruser, ///< Slave ACP - User pins to inform Snoop Control Unit

    // AXI3 Bus Slaves
    axi3_if.slave s_axi_gp0, ///< Slave GP0 - 32-bit data, 32-bit address, 6-bit ID
    axi3_if.slave s_axi_gp1, ///< Slave GP1 - 32-bit data, 32-bit address, 6-bit ID
    axi3_if.slave s_axi_hp0, ///< Slave HP0 - 64-bit data, 32-bit address, 6-bit ID
    axi3_if.slave s_axi_hp1, ///< Slave HP1 - 64-bit data, 32-bit address, 6-bit ID
    axi3_if.slave s_axi_hp2, ///< Slave HP2 - 64-bit data, 32-bit address, 6-bit ID
    axi3_if.slave s_axi_hp3, ///< Slave HP3 - 64-bit data, 32-bit address, 6-bit ID

    // AXI3 Bus Slave FIFO Interfaces
    axi_hp_fifo_if.slave s_axi_hp0_fifo, ///< Slave HP0 - FIFO Control
    axi_hp_fifo_if.slave s_axi_hp1_fifo, ///< Slave HP1 - FIFO Control
    axi_hp_fifo_if.slave s_axi_hp2_fifo, ///< Slave HP2 - FIFO Control
    axi_hp_fifo_if.slave s_axi_hp3_fifo, ///< Slave HP3 - FIFO Control

    // DMA Peripheral Request Interfaces
    dma_req_if.zynq dma0, ///< DMA0 request interface
    dma_req_if.zynq dma1, ///< DMA1 request interface
    dma_req_if.zynq dma2, ///< DMA2 request interface
    dma_req_if.zynq dma3, ///< DMA3 request interface

    // Interrupt Lines
    input  logic [19:0] IRQF2P, ///< Interrupts for processor
    output logic [28:0] IRQP2F, ///< Interrupts for programmable logic

    /// EMIO
    /// Ethernet
    input  logic    eth0_ext_int_in, ///< Ethernet MAC 0 External interrupt
    input  logic    eth1_ext_int_in, ///< Ethernet MAC 1 External interrupt
    gmii_if.mac     eth0,            ///< Ethernet MAC 0 GMII Interface
    gmii_if.mac     eth1,            ///< Ethernet MAC 1 GMII Interface
    ieee1588_if.mac ptp_eth0,        ///< Ethernet MAC 0 PTP output signals
    ieee1588_if.mac ptp_eth1,        ///< Ethernet MAC 1 PTP output signals
    /// JTAG
    jtag.device pjtag, ///< JTAG interface
    /// I2C
    i2c_if.device i2c0, ///< I2C Peripheral 0
    i2c_if.device i2c1, ///< I2C Peripheral 1
    /// SDIO
    sdio_if.master sdio0, ///< SDIO Peripheral 0
    sdio_if.master sdio1, ///< SDIO Peripheral 1
    /// SPI
    spi_if.device spi0, ///< SPI Peripheral 0
    spi_if.device spi1, ///< SPI Peripheral 1
    /// UART
    uart_if.device uart0, ///< UART Peripheral 0
    uart_if.device uart1, ///< UART Peripheral 1
    /// Triple-Timer Counter
    input  logic [2:0] ttc0_CLK, ///< Triple-Timer Counter clock
    output logic [2:0] ttc0_WAVE, ///< Triple-Timer Counter wave output
    input  logic [2:0] ttc1_CLK, ///< Triple-Timer Counter clock
    output logic [2:0] ttc1_WAVE, ///< Triple-Timer Counter wave output
    /// CAN0
    input  logic can0_RX,
    output logic can0_TX,
    /// CAN1
    input  logic can1_RX,
    output logic can1_TX,
    /// GPIO
    input  logic [63:0] gpio_I,
    output logic [63:0] gpio_O,
    output logic [63:0] gpio_TN,
    /// USB0
    output logic [1:0] usb0_PORTINDCTL, ///< Port indicator
    input  logic usb0_VBUSPWRFAULT,     ///< High for USB power fault
    output logic usb0_VBUSPWRSELECT,    ///< Bit to select between system power and external USB power
    /// USB1
    output logic [1:0] usb1_PORTINDCTL, ///< Port indicator
    input  logic usb1_VBUSPWRFAULT,     ///< High for USB power fault
    output logic usb1_VBUSPWRSELECT,    ///< Bit to select between system power and external USB power
    /// WDT - Watchdog Timer
    input  logic wdt_CLKI, ///< Clock input for timer
    output logic wdt_RSTO, ///< Output reset signal

    input  logic sram_int_in, ///< SRAM Interrupt in

    /// Debugging Interfaces
    input  logic [31:0] ftm_debug_f2p, ///< Debugging general-purpose inputs from FPGA
    output logic [31:0] ftm_debug_p2f, ///< Debugging general-purpose outputs to FPGA
    ftm_trigger_if.processor ftm_trigger, ///< Triggers
    ftm_trace_if.processor ftm_trace, ///< Trace logic
    output logic [31:0] trace_DATA, ///< Trace data
    input  logic trace_CLK,         ///< Trace clock
    output logic trace_CTL          ///< Trace control

);

// }}}
///////////////////////////////////////////////////////////////////////////
// Processor Module {{{
///////////////////////////////////////////////////////////////////////////

PS7 processor (
  .DMA0DATYPE(dma0.DATYPE),
  .DMA0DAVALID(dma0.DAVALID),
  .DMA0DRREADY(dma0.DRREADY),
  .DMA0RSTN(dma0.RSTN),
  .DMA1DATYPE(dma1.DATYPE),
  .DMA1DAVALID(dma1.DAVALID),
  .DMA1DRREADY(dma1.DRREADY),
  .DMA1RSTN(dma1.RSTN),
  .DMA2DATYPE(dma2.DATYPE),
  .DMA2DAVALID(dma2.DAVALID),
  .DMA2DRREADY(dma2.DRREADY),
  .DMA2RSTN(dma2.RSTN),
  .DMA3DATYPE(dma3.DATYPE),
  .DMA3DAVALID(dma3.DAVALID),
  .DMA3DRREADY(dma3.DRREADY),
  .DMA3RSTN(dma3.RSTN),
  .EMIOCAN0PHYTX(can0_TX),
  .EMIOCAN1PHYTX(can1_TX),
  .EMIOENET0GMIITXD(eth0.TXD),
  .EMIOENET0GMIITXEN(eth0.TX_EN),
  .EMIOENET0GMIITXER(eth0.TX_ER),
  .EMIOENET0MDIOMDC(eth0.MDIO_MDC),
  .EMIOENET0MDIOO(eth0.MDIO_O),
  .EMIOENET0MDIOTN(eth0.MDIO_TN),
  .EMIOENET0PTPDELAYREQRX(ptp_eth0.DELAYREQRX),
  .EMIOENET0PTPDELAYREQTX(ptp_eth0.DELAYREQTX),
  .EMIOENET0PTPPDELAYREQRX(ptp_eth0.PDELAYREQRX),
  .EMIOENET0PTPPDELAYREQTX(ptp_eth0.PDELAYREQTX),
  .EMIOENET0PTPPDELAYRESPRX(ptp_eth0.PDELAYRESPRX),
  .EMIOENET0PTPPDELAYRESPTX(ptp_eth0.PDELAYRESPTX),
  .EMIOENET0PTPSYNCFRAMERX(ptp_eth0.SYNCFRAMERX),
  .EMIOENET0PTPSYNCFRAMETX(ptp_eth0.SYNCFRAMETX),
  .EMIOENET0SOFRX(ptp_eth0.SOFRX),
  .EMIOENET0SOFTX(ptp_eth0.SOFTX),
  .EMIOENET1GMIITXD(eth1.TXD),
  .EMIOENET1GMIITXEN(eth1.TX_EN),
  .EMIOENET1GMIITXER(eth1.TX_ER),
  .EMIOENET1MDIOMDC(eth1.MDIO_MDC),
  .EMIOENET1MDIOO(eth1.MDIO_O),
  .EMIOENET1MDIOTN(eth1.MDIO_TN),
  .EMIOENET1PTPDELAYREQRX(ptp_eth1.DELAYREQRX),
  .EMIOENET1PTPDELAYREQTX(ptp_eth1.DELAYREQTX),
  .EMIOENET1PTPPDELAYREQRX(ptp_eth1.PDELAYREQRX),
  .EMIOENET1PTPPDELAYREQTX(ptp_eth1.PDELAYREQTX),
  .EMIOENET1PTPPDELAYRESPRX(ptp_eth1.PDELAYRESPRX),
  .EMIOENET1PTPPDELAYRESPTX(ptp_eth1.PDELAYRESPTX),
  .EMIOENET1PTPSYNCFRAMERX(ptp_eth1.SYNCFRAMERX),
  .EMIOENET1PTPSYNCFRAMETX(ptp_eth1.SYNCFRAMETX),
  .EMIOENET1SOFRX(ptp_eth1.SOFRX),
  .EMIOENET1SOFTX(ptp_eth1.SOFTX),
  .EMIOGPIOO(gpio_O),
  .EMIOGPIOTN(gpio_TN),
  .EMIOI2C0SCLO(i2c0.SCLO),
  .EMIOI2C0SCLTN(i2c0.SCLTN),
  .EMIOI2C0SDAO(i2c0.SDAO),
  .EMIOI2C0SDATN(i2c0.SDATN),
  .EMIOI2C1SCLO(i2c1.SCLO),
  .EMIOI2C1SCLTN(i2c1.SCLTN),
  .EMIOI2C1SDAO(i2c1.SDAO),
  .EMIOI2C1SDATN(i2c1.SDATN),
  .EMIOPJTAGTDO(pjtag.TDO),
  .EMIOPJTAGTDTN(pjtag.TDTN),
  .EMIOSDIO0BUSPOW(sdio0.BUSPOW),
  .EMIOSDIO0BUSVOLT(sdio0.BUSVOLT),
  .EMIOSDIO0CLK(sdio0.CLK),
  .EMIOSDIO0CMDO(sdio0.CMDO),
  .EMIOSDIO0CMDTN(sdio0.CMDTN),
  .EMIOSDIO0DATAO(sdio0.DATAO),
  .EMIOSDIO0DATATN(sdio0.DATATN),
  .EMIOSDIO0LED(sdio0.LED),
  .EMIOSDIO1BUSPOW(sdio1.BUSPOW),
  .EMIOSDIO1BUSVOLT(sdio1.BUSVOLT),
  .EMIOSDIO1CLK(sdio1.CLK),
  .EMIOSDIO1CMDO(sdio1.CMDO),
  .EMIOSDIO1CMDTN(sdio1.CMDTN),
  .EMIOSDIO1DATAO(sdio1.DATAO),
  .EMIOSDIO1DATATN(sdio1.DATATN),
  .EMIOSDIO1LED(sdio1.LED),
  .EMIOSPI0MO(spi0.MO),
  .EMIOSPI0MOTN(spi0.MOTN),
  .EMIOSPI0SCLKO(spi0.SCLKO),
  .EMIOSPI0SCLKTN(spi0.SCLKTN),
  .EMIOSPI0SO(spi0.SO),
  .EMIOSPI0SSNTN(spi0.SSNTN),
  .EMIOSPI0SSON(spi0.SSON),
  .EMIOSPI0STN(spi0.STN),
  .EMIOSPI1MO(spi1.MO),
  .EMIOSPI1MOTN(spi1.MOTN),
  .EMIOSPI1SCLKO(spi1.SCLKO),
  .EMIOSPI1SCLKTN(spi1.SCLKTN),
  .EMIOSPI1SO(spi1.SO),
  .EMIOSPI1SSNTN(spi1.SSNTN),
  .EMIOSPI1SSON(spi1.SSON),
  .EMIOSPI1STN(spi1.STN),
  .EMIOTRACECTL(EMIOTRACECTL),
  .EMIOTRACEDATA(EMIOTRACEDATA),
  .EMIOTTC0WAVEO(ttc0_WAVE),
  .EMIOTTC1WAVEO(ttc1_WAVE),
  .EMIOUART0DTRN(uart0.DTRN),
  .EMIOUART0RTSN(uart0.RTSN),
  .EMIOUART0TX(uart0.TX),
  .EMIOUART1DTRN(uart1.DTRN),
  .EMIOUART1RTSN(uart1.RTSN),
  .EMIOUART1TX(uart1.TX),
  .EMIOUSB0PORTINDCTL(EMIOUSB0PORTINDCTL),
  .EMIOUSB0VBUSPWRSELECT(EMIOUSB0VBUSPWRSELECT),
  .EMIOUSB1PORTINDCTL(EMIOUSB1PORTINDCTL),
  .EMIOUSB1VBUSPWRSELECT(EMIOUSB1VBUSPWRSELECT),
  .EMIOWDTRSTO(EMIOWDTRSTO),
  .EVENTEVENTO(EVENTEVENTO),
  .EVENTSTANDBYWFE(EVENTSTANDBYWFE),
  .EVENTSTANDBYWFI(EVENTSTANDBYWFI),
  .FCLKCLK(fclk_CLK),
  .FCLKRESETN(fclk_RESETN),
  .FTMTF2PTRIGACK(ftm_trigger.F2PTRIGACK),
  .FTMTP2FDEBUG(ftm_debug_p2f),
  .FTMTP2FTRIG(ftm_trigger.P2FTRIG),
  .IRQP2F(IRQP2F),
  .MAXIGP0ARADDR(m_axi_gp0.ARADDR),
  .MAXIGP0ARBURST(m_axi_gp0.ARBURST),
  .MAXIGP0ARCACHE(m_axi_gp0.ARCACHE),
  .MAXIGP0ARESETN(m_axi_gp0.ARESETn),
  .MAXIGP0ARID(m_axi_gp0.ARID),
  .MAXIGP0ARLEN(m_axi_gp0.ARLEN),
  .MAXIGP0ARLOCK(m_axi_gp0.ARLOCK),
  .MAXIGP0ARPROT(m_axi_gp0.ARPROT),
  .MAXIGP0ARQOS(m_axi_gp0.ARQOS),
  .MAXIGP0ARSIZE(m_axi_gp0.ARSIZE),
  .MAXIGP0ARVALID(m_axi_gp0.ARVALID),
  .MAXIGP0AWADDR(m_axi_gp0.AWADDR),
  .MAXIGP0AWBURST(m_axi_gp0.AWBURST),
  .MAXIGP0AWCACHE(m_axi_gp0.AWCACHE),
  .MAXIGP0AWID(m_axi_gp0.AWID),
  .MAXIGP0AWLEN(m_axi_gp0.AWLEN),
  .MAXIGP0AWLOCK(m_axi_gp0.AWLOCK),
  .MAXIGP0AWPROT(m_axi_gp0.AWPROT),
  .MAXIGP0AWQOS(m_axi_gp0.AWQOS),
  .MAXIGP0AWSIZE(m_axi_gp0.AWSIZE),
  .MAXIGP0AWVALID(m_axi_gp0.AWVALID),
  .MAXIGP0BREADY(m_axi_gp0.BREADY),
  .MAXIGP0RREADY(m_axi_gp0.RREADY),
  .MAXIGP0WDATA(m_axi_gp0.WDATA),
  .MAXIGP0WID(m_axi_gp0.WID),
  .MAXIGP0WLAST(m_axi_gp0.WLAST),
  .MAXIGP0WSTRB(m_axi_gp0.WSTRB),
  .MAXIGP0WVALID(m_axi_gp0.WVALID),
  .MAXIGP1ARADDR(m_axi_gp1.ARADDR),
  .MAXIGP1ARBURST(m_axi_gp1.ARBURST),
  .MAXIGP1ARCACHE(m_axi_gp1.ARCACHE),
  .MAXIGP1ARESETN(m_axi_gp1.ARESETn),
  .MAXIGP1ARID(m_axi_gp1.ARID),
  .MAXIGP1ARLEN(m_axi_gp1.ARLEN),
  .MAXIGP1ARLOCK(m_axi_gp1.ARLOCK),
  .MAXIGP1ARPROT(m_axi_gp1.ARPROT),
  .MAXIGP1ARQOS(m_axi_gp1.ARQOS),
  .MAXIGP1ARSIZE(m_axi_gp1.ARSIZE),
  .MAXIGP1ARVALID(m_axi_gp1.ARVALID),
  .MAXIGP1AWADDR(m_axi_gp1.AWADDR),
  .MAXIGP1AWBURST(m_axi_gp1.AWBURST),
  .MAXIGP1AWCACHE(m_axi_gp1.AWCACHE),
  .MAXIGP1AWID(m_axi_gp1.AWID),
  .MAXIGP1AWLEN(m_axi_gp1.AWLEN),
  .MAXIGP1AWLOCK(m_axi_gp1.AWLOCK),
  .MAXIGP1AWPROT(m_axi_gp1.AWPROT),
  .MAXIGP1AWQOS(m_axi_gp1.AWQOS),
  .MAXIGP1AWSIZE(m_axi_gp1.AWSIZE),
  .MAXIGP1AWVALID(m_axi_gp1.AWVALID),
  .MAXIGP1BREADY(m_axi_gp1.BREADY),
  .MAXIGP1RREADY(m_axi_gp1.RREADY),
  .MAXIGP1WDATA(m_axi_gp1.WDATA),
  .MAXIGP1WID(m_axi_gp1.WID),
  .MAXIGP1WLAST(m_axi_gp1.WLAST),
  .MAXIGP1WSTRB(m_axi_gp1.WSTRB),
  .MAXIGP1WVALID(m_axi_gp1.WVALID),
  .SAXIACPARESETN(s_axi_acp.ARESETn),
  .SAXIACPARREADY(s_axi_acp.ARREADY),
  .SAXIACPAWREADY(s_axi_acp.AWREADY),
  .SAXIACPBID(s_axi_acp.BID),
  .SAXIACPBRESP(s_axi_acp.BRESP),
  .SAXIACPBVALID(s_axi_acp.BVALID),
  .SAXIACPRDATA(s_axi_acp.RDATA),
  .SAXIACPRID(s_axi_acp.RID),
  .SAXIACPRLAST(s_axi_acp.RLAST),
  .SAXIACPRRESP(s_axi_acp.RRESP),
  .SAXIACPRVALID(s_axi_acp.RVALID),
  .SAXIACPWREADY(s_axi_acp.WREADY),
  .SAXIGP0ARESETN(s_axi_gp0.ARESETn),
  .SAXIGP0ARREADY(s_axi_gp0.ARREADY),
  .SAXIGP0AWREADY(s_axi_gp0.AWREADY),
  .SAXIGP0BID(s_axi_gp0.BID),
  .SAXIGP0BRESP(s_axi_gp0.BRESP),
  .SAXIGP0BVALID(s_axi_gp0.BVALID),
  .SAXIGP0RDATA(s_axi_gp0.RDATA),
  .SAXIGP0RID(s_axi_gp0.RID),
  .SAXIGP0RLAST(s_axi_gp0.RLAST),
  .SAXIGP0RRESP(s_axi_gp0.RRESP),
  .SAXIGP0RVALID(s_axi_gp0.RVALID),
  .SAXIGP0WREADY(s_axi_gp0.WREADY),
  .SAXIGP1ARESETN(s_axi_gp1.ARESETn),
  .SAXIGP1ARREADY(s_axi_gp1.ARREADY),
  .SAXIGP1AWREADY(s_axi_gp1.AWREADY),
  .SAXIGP1BID(s_axi_gp1.BID),
  .SAXIGP1BRESP(s_axi_gp1.BRESP),
  .SAXIGP1BVALID(s_axi_gp1.BVALID),
  .SAXIGP1RDATA(s_axi_gp1.RDATA),
  .SAXIGP1RID(s_axi_gp1.RID),
  .SAXIGP1RLAST(s_axi_gp1.RLAST),
  .SAXIGP1RRESP(s_axi_gp1.RRESP),
  .SAXIGP1RVALID(s_axi_gp1.RVALID),
  .SAXIGP1WREADY(s_axi_gp1.WREADY),
  .SAXIHP0ARESETN(s_axi_hp0.ARESETn),
  .SAXIHP0ARREADY(s_axi_hp0.ARREADY),
  .SAXIHP0AWREADY(s_axi_hp0.AWREADY),
  .SAXIHP0BID(s_axi_hp0.BID),
  .SAXIHP0BRESP(s_axi_hp0.BRESP),
  .SAXIHP0BVALID(s_axi_hp0.BVALID),
  .SAXIHP0RACOUNT(s_axi_hp0_fifo.RACOUNT),
  .SAXIHP0RCOUNT(s_axi_hp0_fifo.RCOUNT),
  .SAXIHP0RDATA(s_axi_hp0.RDATA),
  .SAXIHP0RID(s_axi_hp0.RID),
  .SAXIHP0RLAST(s_axi_hp0.RLAST),
  .SAXIHP0RRESP(s_axi_hp0.RRESP),
  .SAXIHP0RVALID(s_axi_hp0.RVALID),
  .SAXIHP0WACOUNT(s_axi_hp0_fifo.WACOUNT),
  .SAXIHP0WCOUNT(s_axi_hp0_fifo.WCOUNT),
  .SAXIHP0WREADY(s_axi_hp0.WREADY),
  .SAXIHP1ARESETN(s_axi_hp1.ARESETn),
  .SAXIHP1ARREADY(s_axi_hp1.ARREADY),
  .SAXIHP1AWREADY(s_axi_hp1.AWREADY),
  .SAXIHP1BID(s_axi_hp1.BID),
  .SAXIHP1BRESP(s_axi_hp1.BRESP),
  .SAXIHP1BVALID(s_axi_hp1.BVALID),
  .SAXIHP1RACOUNT(s_axi_hp1_fifo.RACOUNT),
  .SAXIHP1RCOUNT(s_axi_hp1_fifo.RCOUNT),
  .SAXIHP1RDATA(s_axi_hp1.RDATA),
  .SAXIHP1RID(s_axi_hp1.RID),
  .SAXIHP1RLAST(s_axi_hp1.RLAST),
  .SAXIHP1RRESP(s_axi_hp1.RRESP),
  .SAXIHP1RVALID(s_axi_hp1.RVALID),
  .SAXIHP1WACOUNT(s_axi_hp1_fifo.WACOUNT),
  .SAXIHP1WCOUNT(s_axi_hp1_fifo.WCOUNT),
  .SAXIHP1WREADY(s_axi_hp1.WREADY),
  .SAXIHP2ARESETN(s_axi_hp2.ARESETn),
  .SAXIHP2ARREADY(s_axi_hp2.ARREADY),
  .SAXIHP2AWREADY(s_axi_hp2.AWREADY),
  .SAXIHP2BID(s_axi_hp2.BID),
  .SAXIHP2BRESP(s_axi_hp2.BRESP),
  .SAXIHP2BVALID(s_axi_hp2.BVALID),
  .SAXIHP2RACOUNT(s_axi_hp2_fifo.RACOUNT),
  .SAXIHP2RCOUNT(s_axi_hp2_fifo.RCOUNT),
  .SAXIHP2RDATA(s_axi_hp2.RDATA),
  .SAXIHP2RID(s_axi_hp2.RID),
  .SAXIHP2RLAST(s_axi_hp2.RLAST),
  .SAXIHP2RRESP(s_axi_hp2.RRESP),
  .SAXIHP2RVALID(s_axi_hp2.RVALID),
  .SAXIHP2WACOUNT(s_axi_hp2_fifo.WACOUNT),
  .SAXIHP2WCOUNT(s_axi_hp2_fifo.WCOUNT),
  .SAXIHP2WREADY(s_axi_hp2.WREADY),
  .SAXIHP3ARESETN(s_axi_hp3.ARESETn),
  .SAXIHP3ARREADY(s_axi_hp3.ARREADY),
  .SAXIHP3AWREADY(s_axi_hp3.AWREADY),
  .SAXIHP3BID(s_axi_hp3.BID),
  .SAXIHP3BRESP(s_axi_hp3.BRESP),
  .SAXIHP3BVALID(s_axi_hp3.BVALID),
  .SAXIHP3RACOUNT(s_axi_hp3_fifo.RACOUNT),
  .SAXIHP3RCOUNT(s_axi_hp3_fifo.RCOUNT),
  .SAXIHP3RDATA(s_axi_hp3.RDATA),
  .SAXIHP3RID(s_axi_hp3.RID),
  .SAXIHP3RLAST(s_axi_hp3.RLAST),
  .SAXIHP3RRESP(s_axi_hp3.RRESP),
  .SAXIHP3RVALID(s_axi_hp3.RVALID),
  .SAXIHP3WACOUNT(s_axi_hp3_fifo.WACOUNT),
  .SAXIHP3WCOUNT(s_axi_hp3_fifo.WCOUNT),
  .SAXIHP3WREADY(s_axi_hp3.WREADY),

  .DDRA(ddr.A),
  .DDRBA(ddr.BA),
  .DDRCASB(ddr.CASB),
  .DDRCKE(ddr.CKE),
  .DDRCKN(ddr.CKN),
  .DDRCKP(ddr.CKP),
  .DDRCSB(ddr.CSB),
  .DDRDM(ddr.DM),
  .DDRDQ(ddr.DQ),
  .DDRDQSN(ddr.DQSN),
  .DDRDQSP(ddr.DQSP),
  .DDRDRSTB(ddr.DRSTB),
  .DDRODT(ddr.ODT),
  .DDRRASB(ddr.RASB),
  .DDRVRN(ddr.VRN),
  .DDRVRP(ddr.VRP),
  .DDRWEB(ddr.WEB),
  .MIO(MIO),
  .PSCLK(PS_CLK),
  .PSPORB(PS_POR_B),
  .PSSRSTB(PS_SRST_B),

  .DDRARB(ddr.ARB),
  .DMA0ACLK(dma0.ACLK),
  .DMA0DAREADY(dma0.DAREADY),
  .DMA0DRLAST(dma0.DRLAST),
  .DMA0DRTYPE(dma0.DRTYPE),
  .DMA0DRVALID(dma0.DRVALID),
  .DMA1ACLK(dma1.ACLK),
  .DMA1DAREADY(dma1.DAREADY),
  .DMA1DRLAST(dma1.DRLAST),
  .DMA1DRTYPE(dma1.DRTYPE),
  .DMA1DRVALID(dma1.DRVALID),
  .DMA2ACLK(dma2.ACLK),
  .DMA2DAREADY(dma2.DAREADY),
  .DMA2DRLAST(dma2.DRLAST),
  .DMA2DRTYPE(dma2.DRTYPE),
  .DMA2DRVALID(dma2.DRVALID),
  .DMA3ACLK(dma3.ACLK),
  .DMA3DAREADY(dma3.DAREADY),
  .DMA3DRLAST(dma3.DRLAST),
  .DMA3DRTYPE(dma3.DRTYPE),
  .DMA3DRVALID(dma3.DRVALID),
  .EMIOCAN0PHYRX(can0_RX),
  .EMIOCAN1PHYRX(can1_RX),
  .EMIOENET0EXTINTIN(eth0_ext_int_in),
  .EMIOENET0GMIICOL(eth0.COL),
  .EMIOENET0GMIICRS(eth0.CRS),
  .EMIOENET0GMIIRXCLK(eth0.RX_CLK),
  .EMIOENET0GMIIRXD(eth0.RXD),
  .EMIOENET0GMIIRXDV(eth0.RX_DV),
  .EMIOENET0GMIIRXER(eth0.RX_ER),
  .EMIOENET0GMIITXCLK(eth0.TX_CLK),
  .EMIOENET0MDIOI(eth0.MDIO_I),
  .EMIOENET1EXTINTIN(eth1_ext_int_in),
  .EMIOENET1GMIICOL(eth1.COL),
  .EMIOENET1GMIICRS(eth1.CRS),
  .EMIOENET1GMIIRXCLK(eth1.RX_CLK),
  .EMIOENET1GMIIRXD(eth1.RXD),
  .EMIOENET1GMIIRXDV(eth1.RX_DV),
  .EMIOENET1GMIIRXER(eth1.RX_ER),
  .EMIOENET1GMIITXCLK(eth1.TX_CLK),
  .EMIOENET1MDIOI(eth1.MDIO_I),
  .EMIOGPIOI(gpio_I),
  .EMIOI2C0SCLI(i2c0.SCLI),
  .EMIOI2C0SDAI(i2c0.SDAI),
  .EMIOI2C1SCLI(i2c1.SCLI),
  .EMIOI2C1SDAI(i2c1.SDAI),
  .EMIOPJTAGTCK(pjtag.TCK),
  .EMIOPJTAGTDI(pjtag.TDI),
  .EMIOPJTAGTMS(pjtag.TMS),
  .EMIOSDIO0CDN(sdio0.CDN),
  .EMIOSDIO0CLKFB(sdio0.CLKFB),
  .EMIOSDIO0CMDI(sdio0.CMDI),
  .EMIOSDIO0DATAI(sdio0.DATAI),
  .EMIOSDIO0WP(sdio0.WP),
  .EMIOSDIO1CDN(sdio1.CDN),
  .EMIOSDIO1CLKFB(sdio1.CLKFB),
  .EMIOSDIO1CMDI(sdio1.CMDI),
  .EMIOSDIO1DATAI(sdio1.DATAI),
  .EMIOSDIO1WP(sdio1.WP),
  .EMIOSPI0MI(spi0.MI),
  .EMIOSPI0SCLKI(spi0.SCLKI),
  .EMIOSPI0SI(spi0.SI),
  .EMIOSPI0SSIN(spi0.SSIN),
  .EMIOSPI1MI(spi1.MI),
  .EMIOSPI1SCLKI(spi1.SCLKI),
  .EMIOSPI1SI(spi1.SI),
  .EMIOSPI1SSIN(spi1.SSIN),
  .EMIOSRAMINTIN(EMIOSRAMINTIN),
  .EMIOTRACECLK(EMIOTRACECLK),
  .EMIOTTC0CLKI(ttc0_CLK),
  .EMIOTTC1CLKI(ttc1_CLK),
  .EMIOUART0CTSN(uart0.CTSN),
  .EMIOUART0DCDN(uart0.DCDN),
  .EMIOUART0DSRN(uart0.DSRN),
  .EMIOUART0RIN(uart0.RIN),
  .EMIOUART0RX(uart0.RX),
  .EMIOUART1CTSN(uart1.CTSN),
  .EMIOUART1DCDN(uart1.DCDN),
  .EMIOUART1DSRN(uart1.DSRN),
  .EMIOUART1RIN(uart1.RIN),
  .EMIOUART1RX(uart1.RX),
  .EMIOUSB0VBUSPWRFAULT(EMIOUSB0VBUSPWRFAULT),
  .EMIOUSB1VBUSPWRFAULT(EMIOUSB1VBUSPWRFAULT),
  .EMIOWDTCLKI(EMIOWDTCLKI),
  .EVENTEVENTI(EVENTEVENTI),
  .FCLKCLKTRIGN(fclk_CLKTRIGN),
  .FPGAIDLEN(FPGAIDLEN),
  .FTMDTRACEINATID(ftm_trace.ATID),
  .FTMDTRACEINCLOCK(ftm_trace.CLOCK),
  .FTMDTRACEINDATA(ftm_trace.DATA),
  .FTMDTRACEINVALID(ftm_trace.VALID),
  .FTMTF2PDEBUG(ftm_debug_f2p),
  .FTMTF2PTRIG(ftm_trigger.F2PTRIG),
  .FTMTP2FTRIGACK(ftm_trigger.P2FTRIGACK),
  .IRQF2P(IRQF2P),
  .MAXIGP0ACLK(m_axi_gp0.ACLK),
  .MAXIGP0ARREADY(m_axi_gp0.ARREADY),
  .MAXIGP0AWREADY(m_axi_gp0.AWREADY),
  .MAXIGP0BID(m_axi_gp0.BID),
  .MAXIGP0BRESP(m_axi_gp0.BRESP),
  .MAXIGP0BVALID(m_axi_gp0.BVALID),
  .MAXIGP0RDATA(m_axi_gp0.RDATA),
  .MAXIGP0RID(m_axi_gp0.RID),
  .MAXIGP0RLAST(m_axi_gp0.RLAST),
  .MAXIGP0RRESP(m_axi_gp0.RRESP),
  .MAXIGP0RVALID(m_axi_gp0.RVALID),
  .MAXIGP0WREADY(m_axi_gp0.WREADY),
  .MAXIGP1ACLK(m_axi_gp1.ACLK),
  .MAXIGP1ARREADY(m_axi_gp1.ARREADY),
  .MAXIGP1AWREADY(m_axi_gp1.AWREADY),
  .MAXIGP1BID(m_axi_gp1.BID),
  .MAXIGP1BRESP(m_axi_gp1.BRESP),
  .MAXIGP1BVALID(m_axi_gp1.BVALID),
  .MAXIGP1RDATA(m_axi_gp1.RDATA),
  .MAXIGP1RID(m_axi_gp1.RID),
  .MAXIGP1RLAST(m_axi_gp1.RLAST),
  .MAXIGP1RRESP(m_axi_gp1.RRESP),
  .MAXIGP1RVALID(m_axi_gp1.RVALID),
  .MAXIGP1WREADY(m_axi_gp1.WREADY),
  .SAXIACPACLK(s_axi_acp.ACLK),
  .SAXIACPARADDR(s_axi_acp.ARADDR),
  .SAXIACPARBURST(s_axi_acp.ARBURST),
  .SAXIACPARCACHE(s_axi_acp.ARCACHE),
  .SAXIACPARID(s_axi_acp.ARID),
  .SAXIACPARLEN(s_axi_acp.ARLEN),
  .SAXIACPARLOCK(s_axi_acp.ARLOCK),
  .SAXIACPARPROT(s_axi_acp.ARPROT),
  .SAXIACPARQOS(s_axi_acp.ARQOS),
  .SAXIACPARSIZE(s_axi_acp.ARSIZE),
  .SAXIACPARUSER(s_axi_acp_aruser),
  .SAXIACPARVALID(s_axi_acp.ARVALID),
  .SAXIACPAWADDR(s_axi_acp.AWADDR),
  .SAXIACPAWBURST(s_axi_acp.AWBURST),
  .SAXIACPAWCACHE(s_axi_acp.AWCACHE),
  .SAXIACPAWID(s_axi_acp.AWID),
  .SAXIACPAWLEN(s_axi_acp.AWLEN),
  .SAXIACPAWLOCK(s_axi_acp.AWLOCK),
  .SAXIACPAWPROT(s_axi_acp.AWPROT),
  .SAXIACPAWQOS(s_axi_acp.AWQOS),
  .SAXIACPAWSIZE(s_axi_acp.AWSIZE),
  .SAXIACPAWUSER(s_axi_acp_awuser),
  .SAXIACPAWVALID(s_axi_acp.AWVALID),
  .SAXIACPBREADY(s_axi_acp.BREADY),
  .SAXIACPRREADY(s_axi_acp.RREADY),
  .SAXIACPWDATA(s_axi_acp.WDATA),
  .SAXIACPWID(s_axi_acp.WID),
  .SAXIACPWLAST(s_axi_acp.WLAST),
  .SAXIACPWSTRB(s_axi_acp.WSTRB),
  .SAXIACPWVALID(s_axi_acp.WVALID),
  .SAXIGP0ACLK(s_axi_gp0.ACLK),
  .SAXIGP0ARADDR(s_axi_gp0.ARADDR),
  .SAXIGP0ARBURST(s_axi_gp0.ARBURST),
  .SAXIGP0ARCACHE(s_axi_gp0.ARCACHE),
  .SAXIGP0ARID(s_axi_gp0.ARID),
  .SAXIGP0ARLEN(s_axi_gp0.ARLEN),
  .SAXIGP0ARLOCK(s_axi_gp0.ARLOCK),
  .SAXIGP0ARPROT(s_axi_gp0.ARPROT),
  .SAXIGP0ARQOS(s_axi_gp0.ARQOS),
  .SAXIGP0ARSIZE(s_axi_gp0.ARSIZE),
  .SAXIGP0ARVALID(s_axi_gp0.ARVALID),
  .SAXIGP0AWADDR(s_axi_gp0.AWADDR),
  .SAXIGP0AWBURST(s_axi_gp0.AWBURST),
  .SAXIGP0AWCACHE(s_axi_gp0.AWCACHE),
  .SAXIGP0AWID(s_axi_gp0.AWID),
  .SAXIGP0AWLEN(s_axi_gp0.AWLEN),
  .SAXIGP0AWLOCK(s_axi_gp0.AWLOCK),
  .SAXIGP0AWPROT(s_axi_gp0.AWPROT),
  .SAXIGP0AWQOS(s_axi_gp0.AWQOS),
  .SAXIGP0AWSIZE(s_axi_gp0.AWSIZE),
  .SAXIGP0AWVALID(s_axi_gp0.AWVALID),
  .SAXIGP0BREADY(s_axi_gp0.BREADY),
  .SAXIGP0RREADY(s_axi_gp0.RREADY),
  .SAXIGP0WDATA(s_axi_gp0.WDATA),
  .SAXIGP0WID(s_axi_gp0.WID),
  .SAXIGP0WLAST(s_axi_gp0.WLAST),
  .SAXIGP0WSTRB(s_axi_gp0.WSTRB),
  .SAXIGP0WVALID(s_axi_gp0.WVALID),
  .SAXIGP1ACLK(s_axi_gp1.ACLK),
  .SAXIGP1ARADDR(s_axi_gp1.ARADDR),
  .SAXIGP1ARBURST(s_axi_gp1.ARBURST),
  .SAXIGP1ARCACHE(s_axi_gp1.ARCACHE),
  .SAXIGP1ARID(s_axi_gp1.ARID),
  .SAXIGP1ARLEN(s_axi_gp1.ARLEN),
  .SAXIGP1ARLOCK(s_axi_gp1.ARLOCK),
  .SAXIGP1ARPROT(s_axi_gp1.ARPROT),
  .SAXIGP1ARQOS(s_axi_gp1.ARQOS),
  .SAXIGP1ARSIZE(s_axi_gp1.ARSIZE),
  .SAXIGP1ARVALID(s_axi_gp1.ARVALID),
  .SAXIGP1AWADDR(s_axi_gp1.AWADDR),
  .SAXIGP1AWBURST(s_axi_gp1.AWBURST),
  .SAXIGP1AWCACHE(s_axi_gp1.AWCACHE),
  .SAXIGP1AWID(s_axi_gp1.AWID),
  .SAXIGP1AWLEN(s_axi_gp1.AWLEN),
  .SAXIGP1AWLOCK(s_axi_gp1.AWLOCK),
  .SAXIGP1AWPROT(s_axi_gp1.AWPROT),
  .SAXIGP1AWQOS(s_axi_gp1.AWQOS),
  .SAXIGP1AWSIZE(s_axi_gp1.AWSIZE),
  .SAXIGP1AWVALID(s_axi_gp1.AWVALID),
  .SAXIGP1BREADY(s_axi_gp1.BREADY),
  .SAXIGP1RREADY(s_axi_gp1.RREADY),
  .SAXIGP1WDATA(s_axi_gp1.WDATA),
  .SAXIGP1WID(s_axi_gp1.WID),
  .SAXIGP1WLAST(s_axi_gp1.WLAST),
  .SAXIGP1WSTRB(s_axi_gp1.WSTRB),
  .SAXIGP1WVALID(s_axi_gp1.WVALID),
  .SAXIHP0ACLK(s_axi_hp0.ACLK),
  .SAXIHP0ARADDR(s_axi_hp0.ARADDR),
  .SAXIHP0ARBURST(s_axi_hp0.ARBURST),
  .SAXIHP0ARCACHE(s_axi_hp0.ARCACHE),
  .SAXIHP0ARID(s_axi_hp0.ARID),
  .SAXIHP0ARLEN(s_axi_hp0.ARLEN),
  .SAXIHP0ARLOCK(s_axi_hp0.ARLOCK),
  .SAXIHP0ARPROT(s_axi_hp0.ARPROT),
  .SAXIHP0ARQOS(s_axi_hp0.ARQOS),
  .SAXIHP0ARSIZE(s_axi_hp0.ARSIZE),
  .SAXIHP0ARVALID(s_axi_hp0.ARVALID),
  .SAXIHP0AWADDR(s_axi_hp0.AWADDR),
  .SAXIHP0AWBURST(s_axi_hp0.AWBURST),
  .SAXIHP0AWCACHE(s_axi_hp0.AWCACHE),
  .SAXIHP0AWID(s_axi_hp0.AWID),
  .SAXIHP0AWLEN(s_axi_hp0.AWLEN),
  .SAXIHP0AWLOCK(s_axi_hp0.AWLOCK),
  .SAXIHP0AWPROT(s_axi_hp0.AWPROT),
  .SAXIHP0AWQOS(s_axi_hp0.AWQOS),
  .SAXIHP0AWSIZE(s_axi_hp0.AWSIZE),
  .SAXIHP0AWVALID(s_axi_hp0.AWVALID),
  .SAXIHP0BREADY(s_axi_hp0.BREADY),
  .SAXIHP0RDISSUECAP1EN(s_axi_hp0_fifo.RDISSUECAP1EN),
  .SAXIHP0RREADY(s_axi_hp0.RREADY),
  .SAXIHP0WDATA(s_axi_hp0.WDATA),
  .SAXIHP0WID(s_axi_hp0.WID),
  .SAXIHP0WLAST(s_axi_hp0.WLAST),
  .SAXIHP0WRISSUECAP1EN(s_axi_hp0_fifo.WRISSUECAP1EN),
  .SAXIHP0WSTRB(s_axi_hp0.WSTRB),
  .SAXIHP0WVALID(s_axi_hp0.WVALID),
  .SAXIHP1ACLK(s_axi_hp1.ACLK),
  .SAXIHP1ARADDR(s_axi_hp1.ARADDR),
  .SAXIHP1ARBURST(s_axi_hp1.ARBURST),
  .SAXIHP1ARCACHE(s_axi_hp1.ARCACHE),
  .SAXIHP1ARID(s_axi_hp1.ARID),
  .SAXIHP1ARLEN(s_axi_hp1.ARLEN),
  .SAXIHP1ARLOCK(s_axi_hp1.ARLOCK),
  .SAXIHP1ARPROT(s_axi_hp1.ARPROT),
  .SAXIHP1ARQOS(s_axi_hp1.ARQOS),
  .SAXIHP1ARSIZE(s_axi_hp1.ARSIZE),
  .SAXIHP1ARVALID(s_axi_hp1.ARVALID),
  .SAXIHP1AWADDR(s_axi_hp1.AWADDR),
  .SAXIHP1AWBURST(s_axi_hp1.AWBURST),
  .SAXIHP1AWCACHE(s_axi_hp1.AWCACHE),
  .SAXIHP1AWID(s_axi_hp1.AWID),
  .SAXIHP1AWLEN(s_axi_hp1.AWLEN),
  .SAXIHP1AWLOCK(s_axi_hp1.AWLOCK),
  .SAXIHP1AWPROT(s_axi_hp1.AWPROT),
  .SAXIHP1AWQOS(s_axi_hp1.AWQOS),
  .SAXIHP1AWSIZE(s_axi_hp1.AWSIZE),
  .SAXIHP1AWVALID(s_axi_hp1.AWVALID),
  .SAXIHP1BREADY(s_axi_hp1.BREADY),
  .SAXIHP1RDISSUECAP1EN(s_axi_hp1_fifo.RDISSUECAP1EN),
  .SAXIHP1RREADY(s_axi_hp1.RREADY),
  .SAXIHP1WDATA(s_axi_hp1.WDATA),
  .SAXIHP1WID(s_axi_hp1.WID),
  .SAXIHP1WLAST(s_axi_hp1.WLAST),
  .SAXIHP1WRISSUECAP1EN(s_axi_hp1_fifo.WRISSUECAP1EN),
  .SAXIHP1WSTRB(s_axi_hp1.WSTRB),
  .SAXIHP1WVALID(s_axi_hp1.WVALID),
  .SAXIHP2ACLK(s_axi_hp2.ACLK),
  .SAXIHP2ARADDR(s_axi_hp2.ARADDR),
  .SAXIHP2ARBURST(s_axi_hp2.ARBURST),
  .SAXIHP2ARCACHE(s_axi_hp2.ARCACHE),
  .SAXIHP2ARID(s_axi_hp2.ARID),
  .SAXIHP2ARLEN(s_axi_hp2.ARLEN),
  .SAXIHP2ARLOCK(s_axi_hp2.ARLOCK),
  .SAXIHP2ARPROT(s_axi_hp2.ARPROT),
  .SAXIHP2ARQOS(s_axi_hp2.ARQOS),
  .SAXIHP2ARSIZE(s_axi_hp2.ARSIZE),
  .SAXIHP2ARVALID(s_axi_hp2.ARVALID),
  .SAXIHP2AWADDR(s_axi_hp2.AWADDR),
  .SAXIHP2AWBURST(s_axi_hp2.AWBURST),
  .SAXIHP2AWCACHE(s_axi_hp2.AWCACHE),
  .SAXIHP2AWID(s_axi_hp2.AWID),
  .SAXIHP2AWLEN(s_axi_hp2.AWLEN),
  .SAXIHP2AWLOCK(s_axi_hp2.AWLOCK),
  .SAXIHP2AWPROT(s_axi_hp2.AWPROT),
  .SAXIHP2AWQOS(s_axi_hp2.AWQOS),
  .SAXIHP2AWSIZE(s_axi_hp2.AWSIZE),
  .SAXIHP2AWVALID(s_axi_hp2.AWVALID),
  .SAXIHP2BREADY(s_axi_hp2.BREADY),
  .SAXIHP2RDISSUECAP1EN(s_axi_hp2_fifo.RDISSUECAP1EN),
  .SAXIHP2RREADY(s_axi_hp2.RREADY),
  .SAXIHP2WDATA(s_axi_hp2.WDATA),
  .SAXIHP2WID(s_axi_hp2.WID),
  .SAXIHP2WLAST(s_axi_hp2.WLAST),
  .SAXIHP2WRISSUECAP1EN(s_axi_hp2_fifo.WRISSUECAP1EN),
  .SAXIHP2WSTRB(s_axi_hp2.WSTRB),
  .SAXIHP2WVALID(s_axi_hp2.WVALID),
  .SAXIHP3ACLK(s_axi_hp3.ACLK),
  .SAXIHP3ARADDR(s_axi_hp3.ARADDR),
  .SAXIHP3ARBURST(s_axi_hp3.ARBURST),
  .SAXIHP3ARCACHE(s_axi_hp3.ARCACHE),
  .SAXIHP3ARID(s_axi_hp3.ARID),
  .SAXIHP3ARLEN(s_axi_hp3.ARLEN),
  .SAXIHP3ARLOCK(s_axi_hp3.ARLOCK),
  .SAXIHP3ARPROT(s_axi_hp3.ARPROT),
  .SAXIHP3ARQOS(s_axi_hp3.ARQOS),
  .SAXIHP3ARSIZE(s_axi_hp3.ARSIZE),
  .SAXIHP3ARVALID(s_axi_hp3.ARVALID),
  .SAXIHP3AWADDR(s_axi_hp3.AWADDR),
  .SAXIHP3AWBURST(s_axi_hp3.AWBURST),
  .SAXIHP3AWCACHE(s_axi_hp3.AWCACHE),
  .SAXIHP3AWID(s_axi_hp3.AWID),
  .SAXIHP3AWLEN(s_axi_hp3.AWLEN),
  .SAXIHP3AWLOCK(s_axi_hp3.AWLOCK),
  .SAXIHP3AWPROT(s_axi_hp3.AWPROT),
  .SAXIHP3AWQOS(s_axi_hp3.AWQOS),
  .SAXIHP3AWSIZE(s_axi_hp3.AWSIZE),
  .SAXIHP3AWVALID(s_axi_hp3.AWVALID),
  .SAXIHP3BREADY(s_axi_hp3.BREADY),
  .SAXIHP3RDISSUECAP1EN(s_axi_hp3_fifo.RDISSUECAP1EN),
  .SAXIHP3RREADY(s_axi_hp3.RREADY),
  .SAXIHP3WDATA(s_axi_hp3.WDATA),
  .SAXIHP3WID(s_axi_hp3.WID),
  .SAXIHP3WLAST(s_axi_hp3.WLAST),
  .SAXIHP3WRISSUECAP1EN(s_axi_hp3_fifo.WRISSUECAP1EN),
  .SAXIHP3WSTRB(s_axi_hp3.WSTRB),
  .SAXIHP3WVALID(s_axi_hp3.WVALID)
);
// }}}

endmodule
/* vim: set fdm=marker: */
