module ps7_wrapper
(
    // AXI3 Bus Masters
    axi3_if.master m_axi_gp0,
    axi3_if.master m_axi_gp1
);

// }}}
///////////////////////////////////////////////////////////////////////////
// Signal Declarations {{{
///////////////////////////////////////////////////////////////////////////

// DDR
wire [31:0] DDRDQ; //inout
wire [14:0] DDRA; //inout
wire [3:0] DDRARB; //input
wire [3:0] DDRDM; //inout
wire [3:0] DDRDQSN; //inout
wire [3:0] DDRDQSP; //inout
wire [2:0] DDRBA; //inout
wire DDRCASB; //inout
wire DDRCKE; //inout
wire DDRCKN; //inout
wire DDRCKP; //inout
wire DDRCSB; //inout
wire DDRDRSTB; //inout
wire DDRODT; //inout
wire DDRRASB; //inout
wire DDRVRN; //inout
wire DDRVRP; //inout
wire DDRWEB; //inout

// DMA0
wire [1:0] DMA0DATYPE; //output
wire [1:0] DMA0DRTYPE; //input
wire DMA0ACLK; //input
wire DMA0DAREADY; //input
wire DMA0DAVALID; //output
wire DMA0DRLAST; //input
wire DMA0DRREADY; //output
wire DMA0DRVALID; //input
wire DMA0RSTN; //output

// DMA1
wire [1:0] DMA1DATYPE; //output
wire [1:0] DMA1DRTYPE; //input
wire DMA1ACLK; //input
wire DMA1DAREADY; //input
wire DMA1DAVALID; //output
wire DMA1DRLAST; //input
wire DMA1DRREADY; //output
wire DMA1DRVALID; //input
wire DMA1RSTN; //output

// DMA2
wire [1:0] DMA2DATYPE; //output
wire [1:0] DMA2DRTYPE; //input
wire DMA2ACLK; //input
wire DMA2DAREADY; //input
wire DMA2DAVALID; //output
wire DMA2DRLAST; //input
wire DMA2DRREADY; //output
wire DMA2DRVALID; //input
wire DMA2RSTN; //output

// DMA3
wire [1:0] DMA3DATYPE; //output
wire [1:0] DMA3DRTYPE; //input
wire DMA3ACLK; //input
wire DMA3DAREADY; //input
wire DMA3DAVALID; //output
wire DMA3DRLAST; //input
wire DMA3DRREADY; //output
wire DMA3DRVALID; //input
wire DMA3RSTN; //output

// EMIOCAN0
wire EMIOCAN0PHYRX; //input
wire EMIOCAN0PHYTX; //output

// EMIOCAN1
wire EMIOCAN1PHYRX; //input
wire EMIOCAN1PHYTX; //output

// EMIOENET0
wire [7:0] EMIOENET0GMIIRXD; //input
wire [7:0] EMIOENET0GMIITXD; //output
wire EMIOENET0EXTINTIN; //input
wire EMIOENET0GMIICOL; //input
wire EMIOENET0GMIICRS; //input
wire EMIOENET0GMIIRXCLK; //input
wire EMIOENET0GMIIRXDV; //input
wire EMIOENET0GMIIRXER; //input
wire EMIOENET0GMIITXCLK; //input
wire EMIOENET0GMIITXEN; //output
wire EMIOENET0GMIITXER; //output
wire EMIOENET0MDIOI; //input
wire EMIOENET0MDIOMDC; //output
wire EMIOENET0MDIOO; //output
wire EMIOENET0MDIOTN; //output
wire EMIOENET0PTPDELAYREQRX; //output
wire EMIOENET0PTPDELAYREQTX; //output
wire EMIOENET0PTPPDELAYREQRX; //output
wire EMIOENET0PTPPDELAYREQTX; //output
wire EMIOENET0PTPPDELAYRESPRX; //output
wire EMIOENET0PTPPDELAYRESPTX; //output
wire EMIOENET0PTPSYNCFRAMERX; //output
wire EMIOENET0PTPSYNCFRAMETX; //output
wire EMIOENET0SOFRX; //output
wire EMIOENET0SOFTX; //output

// EMIOENET1
wire [7:0] EMIOENET1GMIIRXD; //input
wire [7:0] EMIOENET1GMIITXD; //output
wire EMIOENET1EXTINTIN; //input
wire EMIOENET1GMIICOL; //input
wire EMIOENET1GMIICRS; //input
wire EMIOENET1GMIIRXCLK; //input
wire EMIOENET1GMIIRXDV; //input
wire EMIOENET1GMIIRXER; //input
wire EMIOENET1GMIITXCLK; //input
wire EMIOENET1GMIITXEN; //output
wire EMIOENET1GMIITXER; //output
wire EMIOENET1MDIOI; //input
wire EMIOENET1MDIOMDC; //output
wire EMIOENET1MDIOO; //output
wire EMIOENET1MDIOTN; //output
wire EMIOENET1PTPDELAYREQRX; //output
wire EMIOENET1PTPDELAYREQTX; //output
wire EMIOENET1PTPPDELAYREQRX; //output
wire EMIOENET1PTPPDELAYREQTX; //output
wire EMIOENET1PTPPDELAYRESPRX; //output
wire EMIOENET1PTPPDELAYRESPTX; //output
wire EMIOENET1PTPSYNCFRAMERX; //output
wire EMIOENET1PTPSYNCFRAMETX; //output
wire EMIOENET1SOFRX; //output
wire EMIOENET1SOFTX; //output

// EMIOI2C0
wire EMIOI2C0SCLI; //input
wire EMIOI2C0SCLO; //output
wire EMIOI2C0SCLTN; //output
wire EMIOI2C0SDAI; //input
wire EMIOI2C0SDAO; //output
wire EMIOI2C0SDATN; //output

// EMIOI2C1
wire EMIOI2C1SCLI; //input
wire EMIOI2C1SCLO; //output
wire EMIOI2C1SCLTN; //output
wire EMIOI2C1SDAI; //input
wire EMIOI2C1SDAO; //output
wire EMIOI2C1SDATN; //output

// EMIOPJTAG
wire EMIOPJTAGTCK; //input
wire EMIOPJTAGTDI; //input
wire EMIOPJTAGTDO; //output
wire EMIOPJTAGTDTN; //output
wire EMIOPJTAGTMS; //input

// EMIOSDIO0
wire [3:0] EMIOSDIO0DATAI; //input
wire [3:0] EMIOSDIO0DATAO; //output
wire [3:0] EMIOSDIO0DATATN; //output
wire [2:0] EMIOSDIO0BUSVOLT; //output
wire EMIOSDIO0BUSPOW; //output
wire EMIOSDIO0CDN; //input
wire EMIOSDIO0CLK; //output
wire EMIOSDIO0CLKFB; //input
wire EMIOSDIO0CMDI; //input
wire EMIOSDIO0CMDO; //output
wire EMIOSDIO0CMDTN; //output
wire EMIOSDIO0LED; //output
wire EMIOSDIO0WP; //input

// EMIOSDIO1
wire [3:0] EMIOSDIO1DATAI; //input
wire [3:0] EMIOSDIO1DATAO; //output
wire [3:0] EMIOSDIO1DATATN; //output
wire [2:0] EMIOSDIO1BUSVOLT; //output
wire EMIOSDIO1BUSPOW; //output
wire EMIOSDIO1CDN; //input
wire EMIOSDIO1CLK; //output
wire EMIOSDIO1CLKFB; //input
wire EMIOSDIO1CMDI; //input
wire EMIOSDIO1CMDO; //output
wire EMIOSDIO1CMDTN; //output
wire EMIOSDIO1LED; //output
wire EMIOSDIO1WP; //input

// EMIOSPI0
wire [2:0] EMIOSPI0SSON; //output
wire EMIOSPI0MI; //input
wire EMIOSPI0MO; //output
wire EMIOSPI0MOTN; //output
wire EMIOSPI0SCLKI; //input
wire EMIOSPI0SCLKO; //output
wire EMIOSPI0SCLKTN; //output
wire EMIOSPI0SI; //input
wire EMIOSPI0SO; //output
wire EMIOSPI0SSIN; //input
wire EMIOSPI0SSNTN; //output
wire EMIOSPI0STN; //output

// EMIOSPI1
wire [2:0] EMIOSPI1SSON; //output
wire EMIOSPI1MI; //input
wire EMIOSPI1MO; //output
wire EMIOSPI1MOTN; //output
wire EMIOSPI1SCLKI; //input
wire EMIOSPI1SCLKO; //output
wire EMIOSPI1SCLKTN; //output
wire EMIOSPI1SI; //input
wire EMIOSPI1SO; //output
wire EMIOSPI1SSIN; //input
wire EMIOSPI1SSNTN; //output
wire EMIOSPI1STN; //output

// EMIO Misc
wire EMIOSRAMINTIN; //input

// EMIOTRACE
wire [31:0] EMIOTRACEDATA; //output
wire EMIOTRACECLK; //input
wire EMIOTRACECTL; //output

// EMIOUART0
wire EMIOUART0CTSN; //input
wire EMIOUART0DCDN; //input
wire EMIOUART0DSRN; //input
wire EMIOUART0DTRN; //output
wire EMIOUART0RIN; //input
wire EMIOUART0RTSN; //output
wire EMIOUART0RX; //input
wire EMIOUART0TX; //output

// EMIOUART1
wire EMIOUART1CTSN; //input
wire EMIOUART1DCDN; //input
wire EMIOUART1DSRN; //input
wire EMIOUART1DTRN; //output
wire EMIOUART1RIN; //input
wire EMIOUART1RTSN; //output
wire EMIOUART1RX; //input
wire EMIOUART1TX; //output

// EMIOUSB0
wire [1:0] EMIOUSB0PORTINDCTL; //output
wire EMIOUSB0VBUSPWRFAULT; //input
wire EMIOUSB0VBUSPWRSELECT; //output

// EMIOUSB0
wire [1:0] EMIOUSB1PORTINDCTL; //output
wire EMIOUSB1VBUSPWRFAULT; //input
wire EMIOUSB1VBUSPWRSELECT; //output

wire EMIOWDTCLKI; //input
wire EMIOWDTRSTO; //output

// EVENT
wire [1:0] EVENTSTANDBYWFE; //output
wire [1:0] EVENTSTANDBYWFI; //output
wire EVENTEVENTI; //input
wire EVENTEVENTO; //output

wire FPGAIDLEN; //input

// FTM
wire [31:0] FTMDTRACEINDATA; //input
wire [31:0] FTMTF2PDEBUG; //input
wire [31:0] FTMTP2FDEBUG; //output
wire [3:0] FTMDTRACEINATID; //input
wire [3:0] FTMTF2PTRIG; //input
wire [3:0] FTMTF2PTRIGACK; //output
wire [3:0] FTMTP2FTRIG; //output
wire [3:0] FTMTP2FTRIGACK; //input
wire FTMDTRACEINCLOCK; //input
wire FTMDTRACEINVALID; //input

// MAXIGP0
wire [31:0] MAXIGP0ARADDR; //output
wire [31:0] MAXIGP0AWADDR; //output
wire [31:0] MAXIGP0RDATA; //input
wire [31:0] MAXIGP0WDATA; //output
wire [11:0] MAXIGP0ARID; //output
wire [11:0] MAXIGP0AWID; //output
wire [11:0] MAXIGP0BID; //input
wire [11:0] MAXIGP0RID; //input
wire [11:0] MAXIGP0WID; //output
wire [3:0] MAXIGP0ARCACHE; //output
wire [3:0] MAXIGP0ARLEN; //output
wire [3:0] MAXIGP0ARQOS; //output
wire [3:0] MAXIGP0AWCACHE; //output
wire [3:0] MAXIGP0AWLEN; //output
wire [3:0] MAXIGP0AWQOS; //output
wire [3:0] MAXIGP0WSTRB; //output
wire [2:0] MAXIGP0ARPROT; //output
wire [2:0] MAXIGP0AWPROT; //output
wire [1:0] MAXIGP0ARBURST; //output
wire [1:0] MAXIGP0ARLOCK; //output
wire [1:0] MAXIGP0ARSIZE; //output
wire [1:0] MAXIGP0AWBURST; //output
wire [1:0] MAXIGP0AWLOCK; //output
wire [1:0] MAXIGP0AWSIZE; //output
wire [1:0] MAXIGP0BRESP; //input
wire [1:0] MAXIGP0RRESP; //input
wire MAXIGP0ACLK; //input
wire MAXIGP0ARESETN; //output
wire MAXIGP0ARREADY; //input
wire MAXIGP0ARVALID; //output
wire MAXIGP0AWREADY; //input
wire MAXIGP0AWVALID; //output
wire MAXIGP0BREADY; //output
wire MAXIGP0BVALID; //input
wire MAXIGP0RLAST; //input
wire MAXIGP0RREADY; //output
wire MAXIGP0RVALID; //input
wire MAXIGP0WLAST; //output
wire MAXIGP0WREADY; //input
wire MAXIGP0WVALID; //output

// MAXIGP1
wire [31:0] MAXIGP1ARADDR; //output
wire [31:0] MAXIGP1AWADDR; //output
wire [31:0] MAXIGP1RDATA; //input
wire [31:0] MAXIGP1WDATA; //output
wire [11:0] MAXIGP1ARID; //output
wire [11:0] MAXIGP1AWID; //output
wire [11:0] MAXIGP1BID; //input
wire [11:0] MAXIGP1RID; //input
wire [11:0] MAXIGP1WID; //output
wire [3:0] MAXIGP1ARCACHE; //output
wire [3:0] MAXIGP1ARLEN; //output
wire [3:0] MAXIGP1ARQOS; //output
wire [3:0] MAXIGP1AWCACHE; //output
wire [3:0] MAXIGP1AWLEN; //output
wire [3:0] MAXIGP1AWQOS; //output
wire [3:0] MAXIGP1WSTRB; //output
wire [2:0] MAXIGP1ARPROT; //output
wire [2:0] MAXIGP1AWPROT; //output
wire [1:0] MAXIGP1ARBURST; //output
wire [1:0] MAXIGP1ARLOCK; //output
wire [1:0] MAXIGP1ARSIZE; //output
wire [1:0] MAXIGP1AWBURST; //output
wire [1:0] MAXIGP1AWLOCK; //output
wire [1:0] MAXIGP1AWSIZE; //output
wire [1:0] MAXIGP1BRESP; //input
wire [1:0] MAXIGP1RRESP; //input
wire MAXIGP1ACLK; //input
wire MAXIGP1ARESETN; //output
wire MAXIGP1ARREADY; //input
wire MAXIGP1ARVALID; //output
wire MAXIGP1AWREADY; //input
wire MAXIGP1AWVALID; //output
wire MAXIGP1BREADY; //output
wire MAXIGP1BVALID; //input
wire MAXIGP1RLAST; //input
wire MAXIGP1RREADY; //output
wire MAXIGP1RVALID; //input
wire MAXIGP1WLAST; //output
wire MAXIGP1WREADY; //input
wire MAXIGP1WVALID; //output

// PS
wire PSCLK; //inout
wire PSPORB; //inout
wire PSSRSTB; //inout

// SAXIACP
wire [63:0] SAXIACPRDATA; //output
wire [63:0] SAXIACPWDATA; //input
wire [31:0] SAXIACPARADDR; //input
wire [31:0] SAXIACPAWADDR; //input
wire [7:0] SAXIACPWSTRB; //input
wire [3:0] SAXIACPARCACHE; //input
wire [3:0] SAXIACPARLEN; //input
wire [3:0] SAXIACPARQOS; //input
wire [3:0] SAXIACPAWCACHE; //input
wire [3:0] SAXIACPAWLEN; //input
wire [3:0] SAXIACPAWQOS; //input
wire [2:0] SAXIACPARID; //input
wire [2:0] SAXIACPARPROT; //input
wire [2:0] SAXIACPAWID; //input
wire [2:0] SAXIACPAWPROT; //input
wire [2:0] SAXIACPBID; //output
wire [2:0] SAXIACPRID; //output
wire [2:0] SAXIACPWID; //input
wire [1:0] SAXIACPARBURST; //input
wire [1:0] SAXIACPARLOCK; //input
wire [1:0] SAXIACPARSIZE; //input
wire [1:0] SAXIACPAWBURST; //input
wire [1:0] SAXIACPAWLOCK; //input
wire [1:0] SAXIACPAWSIZE; //input
wire [1:0] SAXIACPBRESP; //output
wire [1:0] SAXIACPRRESP; //output
wire SAXIACPACLK; //input
wire SAXIACPARESETN; //output
wire SAXIACPARREADY; //output
wire SAXIACPARVALID; //input
wire SAXIACPAWREADY; //output
wire SAXIACPAWVALID; //input
wire SAXIACPBREADY; //input
wire SAXIACPBVALID; //output
wire SAXIACPRLAST; //output
wire SAXIACPRREADY; //input
wire SAXIACPRVALID; //output
wire SAXIACPWLAST; //input
wire SAXIACPWREADY; //output
wire SAXIACPWVALID; //input

// SAXIGP0
wire [31:0] SAXIGP0ARADDR; //input
wire [31:0] SAXIGP0AWADDR; //input
wire [31:0] SAXIGP0RDATA; //output
wire [31:0] SAXIGP0WDATA; //input
wire [5:0] SAXIGP0ARID; //input
wire [5:0] SAXIGP0AWID; //input
wire [5:0] SAXIGP0BID; //output
wire [5:0] SAXIGP0RID; //output
wire [5:0] SAXIGP0WID; //input
wire [3:0] SAXIGP0ARCACHE; //input
wire [3:0] SAXIGP0ARLEN; //input
wire [3:0] SAXIGP0ARQOS; //input
wire [3:0] SAXIGP0AWCACHE; //input
wire [3:0] SAXIGP0AWLEN; //input
wire [3:0] SAXIGP0AWQOS; //input
wire [3:0] SAXIGP0WSTRB; //input
wire [2:0] SAXIGP0ARPROT; //input
wire [2:0] SAXIGP0AWPROT; //input
wire [1:0] SAXIGP0ARBURST; //input
wire [1:0] SAXIGP0ARLOCK; //input
wire [1:0] SAXIGP0ARSIZE; //input
wire [1:0] SAXIGP0AWBURST; //input
wire [1:0] SAXIGP0AWLOCK; //input
wire [1:0] SAXIGP0AWSIZE; //input
wire [1:0] SAXIGP0BRESP; //output
wire [1:0] SAXIGP0RRESP; //output
wire SAXIGP0ACLK; //input
wire SAXIGP0ARESETN; //output
wire SAXIGP0ARREADY; //output
wire SAXIGP0ARVALID; //input
wire SAXIGP0AWREADY; //output
wire SAXIGP0AWVALID; //input
wire SAXIGP0BREADY; //input
wire SAXIGP0BVALID; //output
wire SAXIGP0RLAST; //output
wire SAXIGP0RREADY; //input
wire SAXIGP0RVALID; //output
wire SAXIGP0WLAST; //input
wire SAXIGP0WREADY; //output
wire SAXIGP0WVALID; //input

// SAXIGP1
wire [31:0] SAXIGP1ARADDR; //input
wire [31:0] SAXIGP1AWADDR; //input
wire [31:0] SAXIGP1RDATA; //output
wire [31:0] SAXIGP1WDATA; //input
wire [5:0] SAXIGP1ARID; //input
wire [5:0] SAXIGP1AWID; //input
wire [5:0] SAXIGP1BID; //output
wire [5:0] SAXIGP1RID; //output
wire [5:0] SAXIGP1WID; //input
wire [3:0] SAXIGP1ARCACHE; //input
wire [3:0] SAXIGP1ARLEN; //input
wire [3:0] SAXIGP1ARQOS; //input
wire [3:0] SAXIGP1AWCACHE; //input
wire [3:0] SAXIGP1AWLEN; //input
wire [3:0] SAXIGP1AWQOS; //input
wire [3:0] SAXIGP1WSTRB; //input
wire [2:0] SAXIGP1ARPROT; //input
wire [2:0] SAXIGP1AWPROT; //input
wire [1:0] SAXIGP1ARBURST; //input
wire [1:0] SAXIGP1ARLOCK; //input
wire [1:0] SAXIGP1ARSIZE; //input
wire [1:0] SAXIGP1AWBURST; //input
wire [1:0] SAXIGP1AWLOCK; //input
wire [1:0] SAXIGP1AWSIZE; //input
wire [1:0] SAXIGP1BRESP; //output
wire [1:0] SAXIGP1RRESP; //output
wire SAXIGP1ACLK; //input
wire SAXIGP1ARESETN; //output
wire SAXIGP1ARREADY; //output
wire SAXIGP1ARVALID; //input
wire SAXIGP1AWREADY; //output
wire SAXIGP1AWVALID; //input
wire SAXIGP1BREADY; //input
wire SAXIGP1BVALID; //output
wire SAXIGP1RLAST; //output
wire SAXIGP1RREADY; //input
wire SAXIGP1RVALID; //output
wire SAXIGP1WLAST; //input
wire SAXIGP1WREADY; //output
wire SAXIGP1WVALID; //input

// SAXIHP0
wire [63:0] SAXIHP0RDATA; //output
wire [63:0] SAXIHP0WDATA; //input
wire [31:0] SAXIHP0ARADDR; //input
wire [31:0] SAXIHP0AWADDR; //input
wire [7:0] SAXIHP0RCOUNT; //output
wire [7:0] SAXIHP0WCOUNT; //output
wire [7:0] SAXIHP0WSTRB; //input
wire [5:0] SAXIHP0ARID; //input
wire [5:0] SAXIHP0AWID; //input
wire [5:0] SAXIHP0BID; //output
wire [5:0] SAXIHP0RID; //output
wire [5:0] SAXIHP0WACOUNT; //output
wire [5:0] SAXIHP0WID; //input
wire [3:0] SAXIHP0ARCACHE; //input
wire [3:0] SAXIHP0ARLEN; //input
wire [3:0] SAXIHP0ARQOS; //input
wire [3:0] SAXIHP0AWCACHE; //input
wire [3:0] SAXIHP0AWLEN; //input
wire [3:0] SAXIHP0AWQOS; //input
wire [2:0] SAXIHP0ARPROT; //input
wire [2:0] SAXIHP0AWPROT; //input
wire [2:0] SAXIHP0RACOUNT; //output
wire [1:0] SAXIHP0ARBURST; //input
wire [1:0] SAXIHP0ARLOCK; //input
wire [1:0] SAXIHP0ARSIZE; //input
wire [1:0] SAXIHP0AWBURST; //input
wire [1:0] SAXIHP0AWLOCK; //input
wire [1:0] SAXIHP0AWSIZE; //input
wire [1:0] SAXIHP0BRESP; //output
wire [1:0] SAXIHP0RRESP; //output
wire SAXIHP0ACLK; //input
wire SAXIHP0ARESETN; //output
wire SAXIHP0ARREADY; //output
wire SAXIHP0ARVALID; //input
wire SAXIHP0AWREADY; //output
wire SAXIHP0AWVALID; //input
wire SAXIHP0BREADY; //input
wire SAXIHP0BVALID; //output
wire SAXIHP0RDISSUECAP1EN; //input
wire SAXIHP0RLAST; //output
wire SAXIHP0RREADY; //input
wire SAXIHP0RVALID; //output
wire SAXIHP0WLAST; //input
wire SAXIHP0WREADY; //output
wire SAXIHP0WRISSUECAP1EN; //input
wire SAXIHP0WVALID; //input

// SAXIHP1
wire [63:0] SAXIHP1RDATA; //output
wire [63:0] SAXIHP1WDATA; //input
wire [31:0] SAXIHP1ARADDR; //input
wire [31:0] SAXIHP1AWADDR; //input
wire [7:0] SAXIHP1RCOUNT; //output
wire [7:0] SAXIHP1WCOUNT; //output
wire [7:0] SAXIHP1WSTRB; //input
wire [5:0] SAXIHP1ARID; //input
wire [5:0] SAXIHP1AWID; //input
wire [5:0] SAXIHP1BID; //output
wire [5:0] SAXIHP1RID; //output
wire [5:0] SAXIHP1WACOUNT; //output
wire [5:0] SAXIHP1WID; //input
wire [3:0] SAXIHP1ARCACHE; //input
wire [3:0] SAXIHP1ARLEN; //input
wire [3:0] SAXIHP1ARQOS; //input
wire [3:0] SAXIHP1AWCACHE; //input
wire [3:0] SAXIHP1AWLEN; //input
wire [3:0] SAXIHP1AWQOS; //input
wire [2:0] SAXIHP1ARPROT; //input
wire [2:0] SAXIHP1AWPROT; //input
wire [2:0] SAXIHP1RACOUNT; //output
wire [1:0] SAXIHP1ARBURST; //input
wire [1:0] SAXIHP1ARLOCK; //input
wire [1:0] SAXIHP1ARSIZE; //input
wire [1:0] SAXIHP1AWBURST; //input
wire [1:0] SAXIHP1AWLOCK; //input
wire [1:0] SAXIHP1AWSIZE; //input
wire [1:0] SAXIHP1BRESP; //output
wire [1:0] SAXIHP1RRESP; //output
wire SAXIHP1ACLK; //input
wire SAXIHP1ARESETN; //output
wire SAXIHP1ARREADY; //output
wire SAXIHP1ARVALID; //input
wire SAXIHP1AWREADY; //output
wire SAXIHP1AWVALID; //input
wire SAXIHP1BREADY; //input
wire SAXIHP1BVALID; //output
wire SAXIHP1RDISSUECAP1EN; //input
wire SAXIHP1RLAST; //output
wire SAXIHP1RREADY; //input
wire SAXIHP1RVALID; //output
wire SAXIHP1WLAST; //input
wire SAXIHP1WREADY; //output
wire SAXIHP1WRISSUECAP1EN; //input
wire SAXIHP1WVALID; //input

// SAXIHP2
wire [63:0] SAXIHP2RDATA; //output
wire [63:0] SAXIHP2WDATA; //input
wire [31:0] SAXIHP2ARADDR; //input
wire [31:0] SAXIHP2AWADDR; //input
wire [7:0] SAXIHP2RCOUNT; //output
wire [7:0] SAXIHP2WCOUNT; //output
wire [7:0] SAXIHP2WSTRB; //input
wire [5:0] SAXIHP2ARID; //input
wire [5:0] SAXIHP2AWID; //input
wire [5:0] SAXIHP2BID; //output
wire [5:0] SAXIHP2RID; //output
wire [5:0] SAXIHP2WACOUNT; //output
wire [5:0] SAXIHP2WID; //input
wire [3:0] SAXIHP2ARCACHE; //input
wire [3:0] SAXIHP2ARLEN; //input
wire [3:0] SAXIHP2ARQOS; //input
wire [3:0] SAXIHP2AWCACHE; //input
wire [3:0] SAXIHP2AWLEN; //input
wire [3:0] SAXIHP2AWQOS; //input
wire [2:0] SAXIHP2ARPROT; //input
wire [2:0] SAXIHP2AWPROT; //input
wire [2:0] SAXIHP2RACOUNT; //output
wire [1:0] SAXIHP2ARBURST; //input
wire [1:0] SAXIHP2ARLOCK; //input
wire [1:0] SAXIHP2ARSIZE; //input
wire [1:0] SAXIHP2AWBURST; //input
wire [1:0] SAXIHP2AWLOCK; //input
wire [1:0] SAXIHP2AWSIZE; //input
wire [1:0] SAXIHP2BRESP; //output
wire [1:0] SAXIHP2RRESP; //output
wire SAXIHP2ACLK; //input
wire SAXIHP2ARESETN; //output
wire SAXIHP2ARREADY; //output
wire SAXIHP2ARVALID; //input
wire SAXIHP2AWREADY; //output
wire SAXIHP2AWVALID; //input
wire SAXIHP2BREADY; //input
wire SAXIHP2BVALID; //output
wire SAXIHP2RDISSUECAP1EN; //input
wire SAXIHP2RLAST; //output
wire SAXIHP2RREADY; //input
wire SAXIHP2RVALID; //output
wire SAXIHP2WLAST; //input
wire SAXIHP2WREADY; //output
wire SAXIHP2WRISSUECAP1EN; //input
wire SAXIHP2WVALID; //input

// SAXIHP3
wire [63:0] SAXIHP3RDATA; //output
wire [63:0] SAXIHP3WDATA; //input
wire [31:0] SAXIHP3ARADDR; //input
wire [31:0] SAXIHP3AWADDR; //input
wire [7:0] SAXIHP3RCOUNT; //output
wire [7:0] SAXIHP3WCOUNT; //output
wire [7:0] SAXIHP3WSTRB; //input
wire [5:0] SAXIHP3ARID; //input
wire [5:0] SAXIHP3AWID; //input
wire [5:0] SAXIHP3BID; //output
wire [5:0] SAXIHP3RID; //output
wire [5:0] SAXIHP3WACOUNT; //output
wire [5:0] SAXIHP3WID; //input
wire [3:0] SAXIHP3ARCACHE; //input
wire [3:0] SAXIHP3ARLEN; //input
wire [3:0] SAXIHP3ARQOS; //input
wire [3:0] SAXIHP3AWCACHE; //input
wire [3:0] SAXIHP3AWLEN; //input
wire [3:0] SAXIHP3AWQOS; //input
wire [2:0] SAXIHP3ARPROT; //input
wire [2:0] SAXIHP3AWPROT; //input
wire [2:0] SAXIHP3RACOUNT; //output
wire [1:0] SAXIHP3ARBURST; //input
wire [1:0] SAXIHP3ARLOCK; //input
wire [1:0] SAXIHP3ARSIZE; //input
wire [1:0] SAXIHP3AWBURST; //input
wire [1:0] SAXIHP3AWLOCK; //input
wire [1:0] SAXIHP3AWSIZE; //input
wire [1:0] SAXIHP3BRESP; //output
wire [1:0] SAXIHP3RRESP; //output
wire SAXIHP3ACLK; //input
wire SAXIHP3ARESETN; //output
wire SAXIHP3ARREADY; //output
wire SAXIHP3ARVALID; //input
wire SAXIHP3AWREADY; //output
wire SAXIHP3AWVALID; //input
wire SAXIHP3BREADY; //input
wire SAXIHP3BVALID; //output
wire SAXIHP3RDISSUECAP1EN; //input
wire SAXIHP3RLAST; //output
wire SAXIHP3RREADY; //input
wire SAXIHP3RVALID; //output
wire SAXIHP3WLAST; //input
wire SAXIHP3WREADY; //output
wire SAXIHP3WRISSUECAP1EN; //input
wire SAXIHP3WVALID; //input

wire [19:0] IRQF2P; //input

wire [28:0] IRQP2F; //output

// EMIOTTC0
wire [2:0] EMIOTTC0CLKI; //input
wire [2:0] EMIOTTC0WAVEO; //output

// EMIOTTC1
wire [2:0] EMIOTTC1CLKI; //input
wire [2:0] EMIOTTC1WAVEO; //output

// FCLK
wire [3:0] FCLKCLK; //output
wire [3:0] FCLKCLKTRIGN; //input
wire [3:0] FCLKRESETN; //output

wire [4:0] SAXIACPARUSER; //input
wire [4:0] SAXIACPAWUSER; //input

wire [53:0] MIO; //inout

// EMIOGPIO
wire [63:0] EMIOGPIOI; //input
wire [63:0] EMIOGPIOO; //output
wire [63:0] EMIOGPIOTN; //output

// }}}
///////////////////////////////////////////////////////////////////////////
// Signal Bundling into Interfaces {{{
///////////////////////////////////////////////////////////////////////////

// MAXIGP0
assign MAXIGP0ACLK = m_axi_gp0.ACLK;
assign MAXIGP0ARESETN = m_axi_gp0.ARESETn;

// Write Address Channel
assign m_axi_gp0.AWID     = MAXIGP0AWID;
assign m_axi_gp0.AWADDR   = MAXIGP0AWADDR;
assign m_axi_gp0.AWLEN    = MAXIGP0AWLEN;
assign m_axi_gp0.AWSIZE   = MAXIGP0AWSIZE;
assign m_axi_gp0.AWBURST  = MAXIGP0AWBURST;
assign m_axi_gp0.AWLOCK   = MAXIGP0AWLOCK;
assign m_axi_gp0.AWCACHE  = MAXIGP0AWCACHE;
assign m_axi_gp0.AWPROT   = MAXIGP0AWPROT;
assign m_axi_gp0.AWVALID  = MAXIGP0AWVALID;
assign MAXIGP0AWREADY     = m_axi_gp0.AWREADY;
// Write Data Channel
assign m_axi_gp0.WID      = MAXIGP0WID;
assign m_axi_gp0.WDATA    = MAXIGP0WDATA;
assign m_axi_gp0.WSTRB    = MAXIGP0WSTRB;
assign m_axi_gp0.WLAST    = MAXIGP0WLAST;
assign m_axi_gp0.WVALID   = MAXIGP0WVALID;
assign MAXIGP0WREADY      = m_axi_gp0.WREADY;
// Write Resposne Channel
assign MAXIGP0BID         = m_axi_gp0.BID;
assign MAXIGP0BRESP       = m_axi_gp0.BRESP;
assign MAXIGP0BVALID      = m_axi_gp0.BVALID;
assign m_axi_gp0.BREADY   = MAXIGP0BREADY;
// Read Address Channel
assign m_axi_gp0.ARID     = MAXIGP0ARID;
assign m_axi_gp0.ARADDR   = MAXIGP0ARADDR;
assign m_axi_gp0.ARLEN    = MAXIGP0ARLEN;
assign m_axi_gp0.ARSIZE   = MAXIGP0ARSIZE;
assign m_axi_gp0.ARBURST  = MAXIGP0ARBURST;
assign m_axi_gp0.ARLOCK   = MAXIGP0ARLOCK;
assign m_axi_gp0.ARCACHE  = MAXIGP0ARCACHE;
assign m_axi_gp0.ARPROT   = MAXIGP0ARPROT;
assign m_axi_gp0.ARVALID  = MAXIGP0ARVALID;
assign MAXIGP0ARREADY     = m_axi_gp0.ARREADY;
// Read Data Channel
assign MAXIGP0RID         = m_axi_gp0.RID;
assign MAXIGP0RDATA       = m_axi_gp0.RDATA;
assign MAXIGP0RRESP       = m_axi_gp0.RRESP;
assign MAXIGP0RLAST       = m_axi_gp0.RLAST;
assign MAXIGP0RVALID      = m_axi_gp0.RVALID;
assign m_axi_gp0.RREADY   = MAXIGP0RREADY;

// MAXIGP1
// Write Address Channel
assign m_axi_gp1.AWID     = MAXIGP1AWID;
assign m_axi_gp1.AWADDR   = MAXIGP1AWADDR;
assign m_axi_gp1.AWLEN    = MAXIGP1AWLEN;
assign m_axi_gp1.AWSIZE   = MAXIGP1AWSIZE;
assign m_axi_gp1.AWBURST  = MAXIGP1AWBURST;
assign m_axi_gp1.AWLOCK   = MAXIGP1AWLOCK;
assign m_axi_gp1.AWCACHE  = MAXIGP1AWCACHE;
assign m_axi_gp1.AWPROT   = MAXIGP1AWPROT;
assign m_axi_gp1.AWVALID  = MAXIGP1AWVALID;
assign MAXIGP1AWREADY     = m_axi_gp1.AWREADY;
// Write Data Channel
assign m_axi_gp1.WID      = MAXIGP1WID;
assign m_axi_gp1.WDATA    = MAXIGP1WDATA;
assign m_axi_gp1.WSTRB    = MAXIGP1WSTRB;
assign m_axi_gp1.WLAST    = MAXIGP1WLAST;
assign m_axi_gp1.WVALID   = MAXIGP1WVALID;
assign MAXIGP1WREADY      = m_axi_gp1.WREADY;
// Write Resposne Channel
assign MAXIGP1BID         = m_axi_gp1.BID;
assign MAXIGP1BRESP       = m_axi_gp1.BRESP;
assign MAXIGP1BVALID      = m_axi_gp1.BVALID;
assign m_axi_gp1.BREADY   = MAXIGP1BREADY;
// Read Address Channel
assign m_axi_gp1.ARID     = MAXIGP1ARID;
assign m_axi_gp1.ARADDR   = MAXIGP1ARADDR;
assign m_axi_gp1.ARLEN    = MAXIGP1ARLEN;
assign m_axi_gp1.ARSIZE   = MAXIGP1ARSIZE;
assign m_axi_gp1.ARBURST  = MAXIGP1ARBURST;
assign m_axi_gp1.ARLOCK   = MAXIGP1ARLOCK;
assign m_axi_gp1.ARCACHE  = MAXIGP1ARCACHE;
assign m_axi_gp1.ARPROT   = MAXIGP1ARPROT;
assign m_axi_gp1.ARVALID  = MAXIGP1ARVALID;
assign MAXIGP1ARREADY     = m_axi_gp1.ARREADY;
// Read Data Channel
assign MAXIGP1RID         = m_axi_gp1.RID;
assign MAXIGP1RDATA       = m_axi_gp1.RDATA;
assign MAXIGP1RRESP       = m_axi_gp1.RRESP;
assign MAXIGP1RLAST       = m_axi_gp1.RLAST;
assign MAXIGP1RVALID      = m_axi_gp1.RVALID;
assign m_axi_gp1.RREADY   = MAXIGP1RREADY;

// }}}
///////////////////////////////////////////////////////////////////////////
// Processor Module {{{
///////////////////////////////////////////////////////////////////////////

PS7 processor (
  .DMA0DATYPE(DMA0DATYPE),
  .DMA0DAVALID(DMA0DAVALID),
  .DMA0DRREADY(DMA0DRREADY),
  .DMA0RSTN(DMA0RSTN),
  .DMA1DATYPE(DMA1DATYPE),
  .DMA1DAVALID(DMA1DAVALID),
  .DMA1DRREADY(DMA1DRREADY),
  .DMA1RSTN(DMA1RSTN),
  .DMA2DATYPE(DMA2DATYPE),
  .DMA2DAVALID(DMA2DAVALID),
  .DMA2DRREADY(DMA2DRREADY),
  .DMA2RSTN(DMA2RSTN),
  .DMA3DATYPE(DMA3DATYPE),
  .DMA3DAVALID(DMA3DAVALID),
  .DMA3DRREADY(DMA3DRREADY),
  .DMA3RSTN(DMA3RSTN),
  .EMIOCAN0PHYTX(EMIOCAN0PHYTX),
  .EMIOCAN1PHYTX(EMIOCAN1PHYTX),
  .EMIOENET0GMIITXD(EMIOENET0GMIITXD),
  .EMIOENET0GMIITXEN(EMIOENET0GMIITXEN),
  .EMIOENET0GMIITXER(EMIOENET0GMIITXER),
  .EMIOENET0MDIOMDC(EMIOENET0MDIOMDC),
  .EMIOENET0MDIOO(EMIOENET0MDIOO),
  .EMIOENET0MDIOTN(EMIOENET0MDIOTN),
  .EMIOENET0PTPDELAYREQRX(EMIOENET0PTPDELAYREQRX),
  .EMIOENET0PTPDELAYREQTX(EMIOENET0PTPDELAYREQTX),
  .EMIOENET0PTPPDELAYREQRX(EMIOENET0PTPPDELAYREQRX),
  .EMIOENET0PTPPDELAYREQTX(EMIOENET0PTPPDELAYREQTX),
  .EMIOENET0PTPPDELAYRESPRX(EMIOENET0PTPPDELAYRESPRX),
  .EMIOENET0PTPPDELAYRESPTX(EMIOENET0PTPPDELAYRESPTX),
  .EMIOENET0PTPSYNCFRAMERX(EMIOENET0PTPSYNCFRAMERX),
  .EMIOENET0PTPSYNCFRAMETX(EMIOENET0PTPSYNCFRAMETX),
  .EMIOENET0SOFRX(EMIOENET0SOFRX),
  .EMIOENET0SOFTX(EMIOENET0SOFTX),
  .EMIOENET1GMIITXD(EMIOENET1GMIITXD),
  .EMIOENET1GMIITXEN(EMIOENET1GMIITXEN),
  .EMIOENET1GMIITXER(EMIOENET1GMIITXER),
  .EMIOENET1MDIOMDC(EMIOENET1MDIOMDC),
  .EMIOENET1MDIOO(EMIOENET1MDIOO),
  .EMIOENET1MDIOTN(EMIOENET1MDIOTN),
  .EMIOENET1PTPDELAYREQRX(EMIOENET1PTPDELAYREQRX),
  .EMIOENET1PTPDELAYREQTX(EMIOENET1PTPDELAYREQTX),
  .EMIOENET1PTPPDELAYREQRX(EMIOENET1PTPPDELAYREQRX),
  .EMIOENET1PTPPDELAYREQTX(EMIOENET1PTPPDELAYREQTX),
  .EMIOENET1PTPPDELAYRESPRX(EMIOENET1PTPPDELAYRESPRX),
  .EMIOENET1PTPPDELAYRESPTX(EMIOENET1PTPPDELAYRESPTX),
  .EMIOENET1PTPSYNCFRAMERX(EMIOENET1PTPSYNCFRAMERX),
  .EMIOENET1PTPSYNCFRAMETX(EMIOENET1PTPSYNCFRAMETX),
  .EMIOENET1SOFRX(EMIOENET1SOFRX),
  .EMIOENET1SOFTX(EMIOENET1SOFTX),
  .EMIOGPIOO(EMIOGPIOO),
  .EMIOGPIOTN(EMIOGPIOTN),
  .EMIOI2C0SCLO(EMIOI2C0SCLO),
  .EMIOI2C0SCLTN(EMIOI2C0SCLTN),
  .EMIOI2C0SDAO(EMIOI2C0SDAO),
  .EMIOI2C0SDATN(EMIOI2C0SDATN),
  .EMIOI2C1SCLO(EMIOI2C1SCLO),
  .EMIOI2C1SCLTN(EMIOI2C1SCLTN),
  .EMIOI2C1SDAO(EMIOI2C1SDAO),
  .EMIOI2C1SDATN(EMIOI2C1SDATN),
  .EMIOPJTAGTDO(EMIOPJTAGTDO),
  .EMIOPJTAGTDTN(EMIOPJTAGTDTN),
  .EMIOSDIO0BUSPOW(EMIOSDIO0BUSPOW),
  .EMIOSDIO0BUSVOLT(EMIOSDIO0BUSVOLT),
  .EMIOSDIO0CLK(EMIOSDIO0CLK),
  .EMIOSDIO0CMDO(EMIOSDIO0CMDO),
  .EMIOSDIO0CMDTN(EMIOSDIO0CMDTN),
  .EMIOSDIO0DATAO(EMIOSDIO0DATAO),
  .EMIOSDIO0DATATN(EMIOSDIO0DATATN),
  .EMIOSDIO0LED(EMIOSDIO0LED),
  .EMIOSDIO1BUSPOW(EMIOSDIO1BUSPOW),
  .EMIOSDIO1BUSVOLT(EMIOSDIO1BUSVOLT),
  .EMIOSDIO1CLK(EMIOSDIO1CLK),
  .EMIOSDIO1CMDO(EMIOSDIO1CMDO),
  .EMIOSDIO1CMDTN(EMIOSDIO1CMDTN),
  .EMIOSDIO1DATAO(EMIOSDIO1DATAO),
  .EMIOSDIO1DATATN(EMIOSDIO1DATATN),
  .EMIOSDIO1LED(EMIOSDIO1LED),
  .EMIOSPI0MO(EMIOSPI0MO),
  .EMIOSPI0MOTN(EMIOSPI0MOTN),
  .EMIOSPI0SCLKO(EMIOSPI0SCLKO),
  .EMIOSPI0SCLKTN(EMIOSPI0SCLKTN),
  .EMIOSPI0SO(EMIOSPI0SO),
  .EMIOSPI0SSNTN(EMIOSPI0SSNTN),
  .EMIOSPI0SSON(EMIOSPI0SSON),
  .EMIOSPI0STN(EMIOSPI0STN),
  .EMIOSPI1MO(EMIOSPI1MO),
  .EMIOSPI1MOTN(EMIOSPI1MOTN),
  .EMIOSPI1SCLKO(EMIOSPI1SCLKO),
  .EMIOSPI1SCLKTN(EMIOSPI1SCLKTN),
  .EMIOSPI1SO(EMIOSPI1SO),
  .EMIOSPI1SSNTN(EMIOSPI1SSNTN),
  .EMIOSPI1SSON(EMIOSPI1SSON),
  .EMIOSPI1STN(EMIOSPI1STN),
  .EMIOTRACECTL(EMIOTRACECTL),
  .EMIOTRACEDATA(EMIOTRACEDATA),
  .EMIOTTC0WAVEO(EMIOTTC0WAVEO),
  .EMIOTTC1WAVEO(EMIOTTC1WAVEO),
  .EMIOUART0DTRN(EMIOUART0DTRN),
  .EMIOUART0RTSN(EMIOUART0RTSN),
  .EMIOUART0TX(EMIOUART0TX),
  .EMIOUART1DTRN(EMIOUART1DTRN),
  .EMIOUART1RTSN(EMIOUART1RTSN),
  .EMIOUART1TX(EMIOUART1TX),
  .EMIOUSB0PORTINDCTL(EMIOUSB0PORTINDCTL),
  .EMIOUSB0VBUSPWRSELECT(EMIOUSB0VBUSPWRSELECT),
  .EMIOUSB1PORTINDCTL(EMIOUSB1PORTINDCTL),
  .EMIOUSB1VBUSPWRSELECT(EMIOUSB1VBUSPWRSELECT),
  .EMIOWDTRSTO(EMIOWDTRSTO),
  .EVENTEVENTO(EVENTEVENTO),
  .EVENTSTANDBYWFE(EVENTSTANDBYWFE),
  .EVENTSTANDBYWFI(EVENTSTANDBYWFI),
  .FCLKCLK(FCLKCLK),
  .FCLKRESETN(FCLKRESETN),
  .FTMTF2PTRIGACK(FTMTF2PTRIGACK),
  .FTMTP2FDEBUG(FTMTP2FDEBUG),
  .FTMTP2FTRIG(FTMTP2FTRIG),
  .IRQP2F(IRQP2F),
  .MAXIGP0ARADDR(MAXIGP0ARADDR),
  .MAXIGP0ARBURST(MAXIGP0ARBURST),
  .MAXIGP0ARCACHE(MAXIGP0ARCACHE),
  .MAXIGP0ARESETN(MAXIGP0ARESETN),
  .MAXIGP0ARID(MAXIGP0ARID),
  .MAXIGP0ARLEN(MAXIGP0ARLEN),
  .MAXIGP0ARLOCK(MAXIGP0ARLOCK),
  .MAXIGP0ARPROT(MAXIGP0ARPROT),
  .MAXIGP0ARQOS(MAXIGP0ARQOS),
  .MAXIGP0ARSIZE(MAXIGP0ARSIZE),
  .MAXIGP0ARVALID(MAXIGP0ARVALID),
  .MAXIGP0AWADDR(MAXIGP0AWADDR),
  .MAXIGP0AWBURST(MAXIGP0AWBURST),
  .MAXIGP0AWCACHE(MAXIGP0AWCACHE),
  .MAXIGP0AWID(MAXIGP0AWID),
  .MAXIGP0AWLEN(MAXIGP0AWLEN),
  .MAXIGP0AWLOCK(MAXIGP0AWLOCK),
  .MAXIGP0AWPROT(MAXIGP0AWPROT),
  .MAXIGP0AWQOS(MAXIGP0AWQOS),
  .MAXIGP0AWSIZE(MAXIGP0AWSIZE),
  .MAXIGP0AWVALID(MAXIGP0AWVALID),
  .MAXIGP0BREADY(MAXIGP0BREADY),
  .MAXIGP0RREADY(MAXIGP0RREADY),
  .MAXIGP0WDATA(MAXIGP0WDATA),
  .MAXIGP0WID(MAXIGP0WID),
  .MAXIGP0WLAST(MAXIGP0WLAST),
  .MAXIGP0WSTRB(MAXIGP0WSTRB),
  .MAXIGP0WVALID(MAXIGP0WVALID),
  .MAXIGP1ARADDR(MAXIGP1ARADDR),
  .MAXIGP1ARBURST(MAXIGP1ARBURST),
  .MAXIGP1ARCACHE(MAXIGP1ARCACHE),
  .MAXIGP1ARESETN(MAXIGP1ARESETN),
  .MAXIGP1ARID(MAXIGP1ARID),
  .MAXIGP1ARLEN(MAXIGP1ARLEN),
  .MAXIGP1ARLOCK(MAXIGP1ARLOCK),
  .MAXIGP1ARPROT(MAXIGP1ARPROT),
  .MAXIGP1ARQOS(MAXIGP1ARQOS),
  .MAXIGP1ARSIZE(MAXIGP1ARSIZE),
  .MAXIGP1ARVALID(MAXIGP1ARVALID),
  .MAXIGP1AWADDR(MAXIGP1AWADDR),
  .MAXIGP1AWBURST(MAXIGP1AWBURST),
  .MAXIGP1AWCACHE(MAXIGP1AWCACHE),
  .MAXIGP1AWID(MAXIGP1AWID),
  .MAXIGP1AWLEN(MAXIGP1AWLEN),
  .MAXIGP1AWLOCK(MAXIGP1AWLOCK),
  .MAXIGP1AWPROT(MAXIGP1AWPROT),
  .MAXIGP1AWQOS(MAXIGP1AWQOS),
  .MAXIGP1AWSIZE(MAXIGP1AWSIZE),
  .MAXIGP1AWVALID(MAXIGP1AWVALID),
  .MAXIGP1BREADY(MAXIGP1BREADY),
  .MAXIGP1RREADY(MAXIGP1RREADY),
  .MAXIGP1WDATA(MAXIGP1WDATA),
  .MAXIGP1WID(MAXIGP1WID),
  .MAXIGP1WLAST(MAXIGP1WLAST),
  .MAXIGP1WSTRB(MAXIGP1WSTRB),
  .MAXIGP1WVALID(MAXIGP1WVALID),
  .SAXIACPARESETN(SAXIACPARESETN),
  .SAXIACPARREADY(SAXIACPARREADY),
  .SAXIACPAWREADY(SAXIACPAWREADY),
  .SAXIACPBID(SAXIACPBID),
  .SAXIACPBRESP(SAXIACPBRESP),
  .SAXIACPBVALID(SAXIACPBVALID),
  .SAXIACPRDATA(SAXIACPRDATA),
  .SAXIACPRID(SAXIACPRID),
  .SAXIACPRLAST(SAXIACPRLAST),
  .SAXIACPRRESP(SAXIACPRRESP),
  .SAXIACPRVALID(SAXIACPRVALID),
  .SAXIACPWREADY(SAXIACPWREADY),
  .SAXIGP0ARESETN(SAXIGP0ARESETN),
  .SAXIGP0ARREADY(SAXIGP0ARREADY),
  .SAXIGP0AWREADY(SAXIGP0AWREADY),
  .SAXIGP0BID(SAXIGP0BID),
  .SAXIGP0BRESP(SAXIGP0BRESP),
  .SAXIGP0BVALID(SAXIGP0BVALID),
  .SAXIGP0RDATA(SAXIGP0RDATA),
  .SAXIGP0RID(SAXIGP0RID),
  .SAXIGP0RLAST(SAXIGP0RLAST),
  .SAXIGP0RRESP(SAXIGP0RRESP),
  .SAXIGP0RVALID(SAXIGP0RVALID),
  .SAXIGP0WREADY(SAXIGP0WREADY),
  .SAXIGP1ARESETN(SAXIGP1ARESETN),
  .SAXIGP1ARREADY(SAXIGP1ARREADY),
  .SAXIGP1AWREADY(SAXIGP1AWREADY),
  .SAXIGP1BID(SAXIGP1BID),
  .SAXIGP1BRESP(SAXIGP1BRESP),
  .SAXIGP1BVALID(SAXIGP1BVALID),
  .SAXIGP1RDATA(SAXIGP1RDATA),
  .SAXIGP1RID(SAXIGP1RID),
  .SAXIGP1RLAST(SAXIGP1RLAST),
  .SAXIGP1RRESP(SAXIGP1RRESP),
  .SAXIGP1RVALID(SAXIGP1RVALID),
  .SAXIGP1WREADY(SAXIGP1WREADY),
  .SAXIHP0ARESETN(SAXIHP0ARESETN),
  .SAXIHP0ARREADY(SAXIHP0ARREADY),
  .SAXIHP0AWREADY(SAXIHP0AWREADY),
  .SAXIHP0BID(SAXIHP0BID),
  .SAXIHP0BRESP(SAXIHP0BRESP),
  .SAXIHP0BVALID(SAXIHP0BVALID),
  .SAXIHP0RACOUNT(SAXIHP0RACOUNT),
  .SAXIHP0RCOUNT(SAXIHP0RCOUNT),
  .SAXIHP0RDATA(SAXIHP0RDATA),
  .SAXIHP0RID(SAXIHP0RID),
  .SAXIHP0RLAST(SAXIHP0RLAST),
  .SAXIHP0RRESP(SAXIHP0RRESP),
  .SAXIHP0RVALID(SAXIHP0RVALID),
  .SAXIHP0WACOUNT(SAXIHP0WACOUNT),
  .SAXIHP0WCOUNT(SAXIHP0WCOUNT),
  .SAXIHP0WREADY(SAXIHP0WREADY),
  .SAXIHP1ARESETN(SAXIHP1ARESETN),
  .SAXIHP1ARREADY(SAXIHP1ARREADY),
  .SAXIHP1AWREADY(SAXIHP1AWREADY),
  .SAXIHP1BID(SAXIHP1BID),
  .SAXIHP1BRESP(SAXIHP1BRESP),
  .SAXIHP1BVALID(SAXIHP1BVALID),
  .SAXIHP1RACOUNT(SAXIHP1RACOUNT),
  .SAXIHP1RCOUNT(SAXIHP1RCOUNT),
  .SAXIHP1RDATA(SAXIHP1RDATA),
  .SAXIHP1RID(SAXIHP1RID),
  .SAXIHP1RLAST(SAXIHP1RLAST),
  .SAXIHP1RRESP(SAXIHP1RRESP),
  .SAXIHP1RVALID(SAXIHP1RVALID),
  .SAXIHP1WACOUNT(SAXIHP1WACOUNT),
  .SAXIHP1WCOUNT(SAXIHP1WCOUNT),
  .SAXIHP1WREADY(SAXIHP1WREADY),
  .SAXIHP2ARESETN(SAXIHP2ARESETN),
  .SAXIHP2ARREADY(SAXIHP2ARREADY),
  .SAXIHP2AWREADY(SAXIHP2AWREADY),
  .SAXIHP2BID(SAXIHP2BID),
  .SAXIHP2BRESP(SAXIHP2BRESP),
  .SAXIHP2BVALID(SAXIHP2BVALID),
  .SAXIHP2RACOUNT(SAXIHP2RACOUNT),
  .SAXIHP2RCOUNT(SAXIHP2RCOUNT),
  .SAXIHP2RDATA(SAXIHP2RDATA),
  .SAXIHP2RID(SAXIHP2RID),
  .SAXIHP2RLAST(SAXIHP2RLAST),
  .SAXIHP2RRESP(SAXIHP2RRESP),
  .SAXIHP2RVALID(SAXIHP2RVALID),
  .SAXIHP2WACOUNT(SAXIHP2WACOUNT),
  .SAXIHP2WCOUNT(SAXIHP2WCOUNT),
  .SAXIHP2WREADY(SAXIHP2WREADY),
  .SAXIHP3ARESETN(SAXIHP3ARESETN),
  .SAXIHP3ARREADY(SAXIHP3ARREADY),
  .SAXIHP3AWREADY(SAXIHP3AWREADY),
  .SAXIHP3BID(SAXIHP3BID),
  .SAXIHP3BRESP(SAXIHP3BRESP),
  .SAXIHP3BVALID(SAXIHP3BVALID),
  .SAXIHP3RACOUNT(SAXIHP3RACOUNT),
  .SAXIHP3RCOUNT(SAXIHP3RCOUNT),
  .SAXIHP3RDATA(SAXIHP3RDATA),
  .SAXIHP3RID(SAXIHP3RID),
  .SAXIHP3RLAST(SAXIHP3RLAST),
  .SAXIHP3RRESP(SAXIHP3RRESP),
  .SAXIHP3RVALID(SAXIHP3RVALID),
  .SAXIHP3WACOUNT(SAXIHP3WACOUNT),
  .SAXIHP3WCOUNT(SAXIHP3WCOUNT),
  .SAXIHP3WREADY(SAXIHP3WREADY),

  .DDRA(DDRA),
  .DDRBA(DDRBA),
  .DDRCASB(DDRCASB),
  .DDRCKE(DDRCKE),
  .DDRCKN(DDRCKN),
  .DDRCKP(DDRCKP),
  .DDRCSB(DDRCSB),
  .DDRDM(DDRDM),
  .DDRDQ(DDRDQ),
  .DDRDQSN(DDRDQSN),
  .DDRDQSP(DDRDQSP),
  .DDRDRSTB(DDRDRSTB),
  .DDRODT(DDRODT),
  .DDRRASB(DDRRASB),
  .DDRVRN(DDRVRN),
  .DDRVRP(DDRVRP),
  .DDRWEB(DDRWEB),
  .MIO(MIO),
  .PSCLK(PSCLK),
  .PSPORB(PSPORB),
  .PSSRSTB(PSSRSTB),

  .DDRARB(DDRARB),
  .DMA0ACLK(DMA0ACLK),
  .DMA0DAREADY(DMA0DAREADY),
  .DMA0DRLAST(DMA0DRLAST),
  .DMA0DRTYPE(DMA0DRTYPE),
  .DMA0DRVALID(DMA0DRVALID),
  .DMA1ACLK(DMA1ACLK),
  .DMA1DAREADY(DMA1DAREADY),
  .DMA1DRLAST(DMA1DRLAST),
  .DMA1DRTYPE(DMA1DRTYPE),
  .DMA1DRVALID(DMA1DRVALID),
  .DMA2ACLK(DMA2ACLK),
  .DMA2DAREADY(DMA2DAREADY),
  .DMA2DRLAST(DMA2DRLAST),
  .DMA2DRTYPE(DMA2DRTYPE),
  .DMA2DRVALID(DMA2DRVALID),
  .DMA3ACLK(DMA3ACLK),
  .DMA3DAREADY(DMA3DAREADY),
  .DMA3DRLAST(DMA3DRLAST),
  .DMA3DRTYPE(DMA3DRTYPE),
  .DMA3DRVALID(DMA3DRVALID),
  .EMIOCAN0PHYRX(EMIOCAN0PHYRX),
  .EMIOCAN1PHYRX(EMIOCAN1PHYRX),
  .EMIOENET0EXTINTIN(EMIOENET0EXTINTIN),
  .EMIOENET0GMIICOL(EMIOENET0GMIICOL),
  .EMIOENET0GMIICRS(EMIOENET0GMIICRS),
  .EMIOENET0GMIIRXCLK(EMIOENET0GMIIRXCLK),
  .EMIOENET0GMIIRXD(EMIOENET0GMIIRXD),
  .EMIOENET0GMIIRXDV(EMIOENET0GMIIRXDV),
  .EMIOENET0GMIIRXER(EMIOENET0GMIIRXER),
  .EMIOENET0GMIITXCLK(EMIOENET0GMIITXCLK),
  .EMIOENET0MDIOI(EMIOENET0MDIOI),
  .EMIOENET1EXTINTIN(EMIOENET1EXTINTIN),
  .EMIOENET1GMIICOL(EMIOENET1GMIICOL),
  .EMIOENET1GMIICRS(EMIOENET1GMIICRS),
  .EMIOENET1GMIIRXCLK(EMIOENET1GMIIRXCLK),
  .EMIOENET1GMIIRXD(EMIOENET1GMIIRXD),
  .EMIOENET1GMIIRXDV(EMIOENET1GMIIRXDV),
  .EMIOENET1GMIIRXER(EMIOENET1GMIIRXER),
  .EMIOENET1GMIITXCLK(EMIOENET1GMIITXCLK),
  .EMIOENET1MDIOI(EMIOENET1MDIOI),
  .EMIOGPIOI(EMIOGPIOI),
  .EMIOI2C0SCLI(EMIOI2C0SCLI),
  .EMIOI2C0SDAI(EMIOI2C0SDAI),
  .EMIOI2C1SCLI(EMIOI2C1SCLI),
  .EMIOI2C1SDAI(EMIOI2C1SDAI),
  .EMIOPJTAGTCK(EMIOPJTAGTCK),
  .EMIOPJTAGTDI(EMIOPJTAGTDI),
  .EMIOPJTAGTMS(EMIOPJTAGTMS),
  .EMIOSDIO0CDN(EMIOSDIO0CDN),
  .EMIOSDIO0CLKFB(EMIOSDIO0CLKFB),
  .EMIOSDIO0CMDI(EMIOSDIO0CMDI),
  .EMIOSDIO0DATAI(EMIOSDIO0DATAI),
  .EMIOSDIO0WP(EMIOSDIO0WP),
  .EMIOSDIO1CDN(EMIOSDIO1CDN),
  .EMIOSDIO1CLKFB(EMIOSDIO1CLKFB),
  .EMIOSDIO1CMDI(EMIOSDIO1CMDI),
  .EMIOSDIO1DATAI(EMIOSDIO1DATAI),
  .EMIOSDIO1WP(EMIOSDIO1WP),
  .EMIOSPI0MI(EMIOSPI0MI),
  .EMIOSPI0SCLKI(EMIOSPI0SCLKI),
  .EMIOSPI0SI(EMIOSPI0SI),
  .EMIOSPI0SSIN(EMIOSPI0SSIN),
  .EMIOSPI1MI(EMIOSPI1MI),
  .EMIOSPI1SCLKI(EMIOSPI1SCLKI),
  .EMIOSPI1SI(EMIOSPI1SI),
  .EMIOSPI1SSIN(EMIOSPI1SSIN),
  .EMIOSRAMINTIN(EMIOSRAMINTIN),
  .EMIOTRACECLK(EMIOTRACECLK),
  .EMIOTTC0CLKI(EMIOTTC0CLKI),
  .EMIOTTC1CLKI(EMIOTTC1CLKI),
  .EMIOUART0CTSN(EMIOUART0CTSN),
  .EMIOUART0DCDN(EMIOUART0DCDN),
  .EMIOUART0DSRN(EMIOUART0DSRN),
  .EMIOUART0RIN(EMIOUART0RIN),
  .EMIOUART0RX(EMIOUART0RX),
  .EMIOUART1CTSN(EMIOUART1CTSN),
  .EMIOUART1DCDN(EMIOUART1DCDN),
  .EMIOUART1DSRN(EMIOUART1DSRN),
  .EMIOUART1RIN(EMIOUART1RIN),
  .EMIOUART1RX(EMIOUART1RX),
  .EMIOUSB0VBUSPWRFAULT(EMIOUSB0VBUSPWRFAULT),
  .EMIOUSB1VBUSPWRFAULT(EMIOUSB1VBUSPWRFAULT),
  .EMIOWDTCLKI(EMIOWDTCLKI),
  .EVENTEVENTI(EVENTEVENTI),
  .FCLKCLKTRIGN(FCLKCLKTRIGN),
  .FPGAIDLEN(FPGAIDLEN),
  .FTMDTRACEINATID(FTMDTRACEINATID),
  .FTMDTRACEINCLOCK(FTMDTRACEINCLOCK),
  .FTMDTRACEINDATA(FTMDTRACEINDATA),
  .FTMDTRACEINVALID(FTMDTRACEINVALID),
  .FTMTF2PDEBUG(FTMTF2PDEBUG),
  .FTMTF2PTRIG(FTMTF2PTRIG),
  .FTMTP2FTRIGACK(FTMTP2FTRIGACK),
  .IRQF2P(IRQF2P),
  .MAXIGP0ACLK(MAXIGP0ACLK),
  .MAXIGP0ARREADY(MAXIGP0ARREADY),
  .MAXIGP0AWREADY(MAXIGP0AWREADY),
  .MAXIGP0BID(MAXIGP0BID),
  .MAXIGP0BRESP(MAXIGP0BRESP),
  .MAXIGP0BVALID(MAXIGP0BVALID),
  .MAXIGP0RDATA(MAXIGP0RDATA),
  .MAXIGP0RID(MAXIGP0RID),
  .MAXIGP0RLAST(MAXIGP0RLAST),
  .MAXIGP0RRESP(MAXIGP0RRESP),
  .MAXIGP0RVALID(MAXIGP0RVALID),
  .MAXIGP0WREADY(MAXIGP0WREADY),
  .MAXIGP1ACLK(MAXIGP1ACLK),
  .MAXIGP1ARREADY(MAXIGP1ARREADY),
  .MAXIGP1AWREADY(MAXIGP1AWREADY),
  .MAXIGP1BID(MAXIGP1BID),
  .MAXIGP1BRESP(MAXIGP1BRESP),
  .MAXIGP1BVALID(MAXIGP1BVALID),
  .MAXIGP1RDATA(MAXIGP1RDATA),
  .MAXIGP1RID(MAXIGP1RID),
  .MAXIGP1RLAST(MAXIGP1RLAST),
  .MAXIGP1RRESP(MAXIGP1RRESP),
  .MAXIGP1RVALID(MAXIGP1RVALID),
  .MAXIGP1WREADY(MAXIGP1WREADY),
  .SAXIACPACLK(SAXIACPACLK),
  .SAXIACPARADDR(SAXIACPARADDR),
  .SAXIACPARBURST(SAXIACPARBURST),
  .SAXIACPARCACHE(SAXIACPARCACHE),
  .SAXIACPARID(SAXIACPARID),
  .SAXIACPARLEN(SAXIACPARLEN),
  .SAXIACPARLOCK(SAXIACPARLOCK),
  .SAXIACPARPROT(SAXIACPARPROT),
  .SAXIACPARQOS(SAXIACPARQOS),
  .SAXIACPARSIZE(SAXIACPARSIZE),
  .SAXIACPARUSER(SAXIACPARUSER),
  .SAXIACPARVALID(SAXIACPARVALID),
  .SAXIACPAWADDR(SAXIACPAWADDR),
  .SAXIACPAWBURST(SAXIACPAWBURST),
  .SAXIACPAWCACHE(SAXIACPAWCACHE),
  .SAXIACPAWID(SAXIACPAWID),
  .SAXIACPAWLEN(SAXIACPAWLEN),
  .SAXIACPAWLOCK(SAXIACPAWLOCK),
  .SAXIACPAWPROT(SAXIACPAWPROT),
  .SAXIACPAWQOS(SAXIACPAWQOS),
  .SAXIACPAWSIZE(SAXIACPAWSIZE),
  .SAXIACPAWUSER(SAXIACPAWUSER),
  .SAXIACPAWVALID(SAXIACPAWVALID),
  .SAXIACPBREADY(SAXIACPBREADY),
  .SAXIACPRREADY(SAXIACPRREADY),
  .SAXIACPWDATA(SAXIACPWDATA),
  .SAXIACPWID(SAXIACPWID),
  .SAXIACPWLAST(SAXIACPWLAST),
  .SAXIACPWSTRB(SAXIACPWSTRB),
  .SAXIACPWVALID(SAXIACPWVALID),
  .SAXIGP0ACLK(SAXIGP0ACLK),
  .SAXIGP0ARADDR(SAXIGP0ARADDR),
  .SAXIGP0ARBURST(SAXIGP0ARBURST),
  .SAXIGP0ARCACHE(SAXIGP0ARCACHE),
  .SAXIGP0ARID(SAXIGP0ARID),
  .SAXIGP0ARLEN(SAXIGP0ARLEN),
  .SAXIGP0ARLOCK(SAXIGP0ARLOCK),
  .SAXIGP0ARPROT(SAXIGP0ARPROT),
  .SAXIGP0ARQOS(SAXIGP0ARQOS),
  .SAXIGP0ARSIZE(SAXIGP0ARSIZE),
  .SAXIGP0ARVALID(SAXIGP0ARVALID),
  .SAXIGP0AWADDR(SAXIGP0AWADDR),
  .SAXIGP0AWBURST(SAXIGP0AWBURST),
  .SAXIGP0AWCACHE(SAXIGP0AWCACHE),
  .SAXIGP0AWID(SAXIGP0AWID),
  .SAXIGP0AWLEN(SAXIGP0AWLEN),
  .SAXIGP0AWLOCK(SAXIGP0AWLOCK),
  .SAXIGP0AWPROT(SAXIGP0AWPROT),
  .SAXIGP0AWQOS(SAXIGP0AWQOS),
  .SAXIGP0AWSIZE(SAXIGP0AWSIZE),
  .SAXIGP0AWVALID(SAXIGP0AWVALID),
  .SAXIGP0BREADY(SAXIGP0BREADY),
  .SAXIGP0RREADY(SAXIGP0RREADY),
  .SAXIGP0WDATA(SAXIGP0WDATA),
  .SAXIGP0WID(SAXIGP0WID),
  .SAXIGP0WLAST(SAXIGP0WLAST),
  .SAXIGP0WSTRB(SAXIGP0WSTRB),
  .SAXIGP0WVALID(SAXIGP0WVALID),
  .SAXIGP1ACLK(SAXIGP1ACLK),
  .SAXIGP1ARADDR(SAXIGP1ARADDR),
  .SAXIGP1ARBURST(SAXIGP1ARBURST),
  .SAXIGP1ARCACHE(SAXIGP1ARCACHE),
  .SAXIGP1ARID(SAXIGP1ARID),
  .SAXIGP1ARLEN(SAXIGP1ARLEN),
  .SAXIGP1ARLOCK(SAXIGP1ARLOCK),
  .SAXIGP1ARPROT(SAXIGP1ARPROT),
  .SAXIGP1ARQOS(SAXIGP1ARQOS),
  .SAXIGP1ARSIZE(SAXIGP1ARSIZE),
  .SAXIGP1ARVALID(SAXIGP1ARVALID),
  .SAXIGP1AWADDR(SAXIGP1AWADDR),
  .SAXIGP1AWBURST(SAXIGP1AWBURST),
  .SAXIGP1AWCACHE(SAXIGP1AWCACHE),
  .SAXIGP1AWID(SAXIGP1AWID),
  .SAXIGP1AWLEN(SAXIGP1AWLEN),
  .SAXIGP1AWLOCK(SAXIGP1AWLOCK),
  .SAXIGP1AWPROT(SAXIGP1AWPROT),
  .SAXIGP1AWQOS(SAXIGP1AWQOS),
  .SAXIGP1AWSIZE(SAXIGP1AWSIZE),
  .SAXIGP1AWVALID(SAXIGP1AWVALID),
  .SAXIGP1BREADY(SAXIGP1BREADY),
  .SAXIGP1RREADY(SAXIGP1RREADY),
  .SAXIGP1WDATA(SAXIGP1WDATA),
  .SAXIGP1WID(SAXIGP1WID),
  .SAXIGP1WLAST(SAXIGP1WLAST),
  .SAXIGP1WSTRB(SAXIGP1WSTRB),
  .SAXIGP1WVALID(SAXIGP1WVALID),
  .SAXIHP0ACLK(SAXIHP0ACLK),
  .SAXIHP0ARADDR(SAXIHP0ARADDR),
  .SAXIHP0ARBURST(SAXIHP0ARBURST),
  .SAXIHP0ARCACHE(SAXIHP0ARCACHE),
  .SAXIHP0ARID(SAXIHP0ARID),
  .SAXIHP0ARLEN(SAXIHP0ARLEN),
  .SAXIHP0ARLOCK(SAXIHP0ARLOCK),
  .SAXIHP0ARPROT(SAXIHP0ARPROT),
  .SAXIHP0ARQOS(SAXIHP0ARQOS),
  .SAXIHP0ARSIZE(SAXIHP0ARSIZE),
  .SAXIHP0ARVALID(SAXIHP0ARVALID),
  .SAXIHP0AWADDR(SAXIHP0AWADDR),
  .SAXIHP0AWBURST(SAXIHP0AWBURST),
  .SAXIHP0AWCACHE(SAXIHP0AWCACHE),
  .SAXIHP0AWID(SAXIHP0AWID),
  .SAXIHP0AWLEN(SAXIHP0AWLEN),
  .SAXIHP0AWLOCK(SAXIHP0AWLOCK),
  .SAXIHP0AWPROT(SAXIHP0AWPROT),
  .SAXIHP0AWQOS(SAXIHP0AWQOS),
  .SAXIHP0AWSIZE(SAXIHP0AWSIZE),
  .SAXIHP0AWVALID(SAXIHP0AWVALID),
  .SAXIHP0BREADY(SAXIHP0BREADY),
  .SAXIHP0RDISSUECAP1EN(SAXIHP0RDISSUECAP1EN),
  .SAXIHP0RREADY(SAXIHP0RREADY),
  .SAXIHP0WDATA(SAXIHP0WDATA),
  .SAXIHP0WID(SAXIHP0WID),
  .SAXIHP0WLAST(SAXIHP0WLAST),
  .SAXIHP0WRISSUECAP1EN(SAXIHP0WRISSUECAP1EN),
  .SAXIHP0WSTRB(SAXIHP0WSTRB),
  .SAXIHP0WVALID(SAXIHP0WVALID),
  .SAXIHP1ACLK(SAXIHP1ACLK),
  .SAXIHP1ARADDR(SAXIHP1ARADDR),
  .SAXIHP1ARBURST(SAXIHP1ARBURST),
  .SAXIHP1ARCACHE(SAXIHP1ARCACHE),
  .SAXIHP1ARID(SAXIHP1ARID),
  .SAXIHP1ARLEN(SAXIHP1ARLEN),
  .SAXIHP1ARLOCK(SAXIHP1ARLOCK),
  .SAXIHP1ARPROT(SAXIHP1ARPROT),
  .SAXIHP1ARQOS(SAXIHP1ARQOS),
  .SAXIHP1ARSIZE(SAXIHP1ARSIZE),
  .SAXIHP1ARVALID(SAXIHP1ARVALID),
  .SAXIHP1AWADDR(SAXIHP1AWADDR),
  .SAXIHP1AWBURST(SAXIHP1AWBURST),
  .SAXIHP1AWCACHE(SAXIHP1AWCACHE),
  .SAXIHP1AWID(SAXIHP1AWID),
  .SAXIHP1AWLEN(SAXIHP1AWLEN),
  .SAXIHP1AWLOCK(SAXIHP1AWLOCK),
  .SAXIHP1AWPROT(SAXIHP1AWPROT),
  .SAXIHP1AWQOS(SAXIHP1AWQOS),
  .SAXIHP1AWSIZE(SAXIHP1AWSIZE),
  .SAXIHP1AWVALID(SAXIHP1AWVALID),
  .SAXIHP1BREADY(SAXIHP1BREADY),
  .SAXIHP1RDISSUECAP1EN(SAXIHP1RDISSUECAP1EN),
  .SAXIHP1RREADY(SAXIHP1RREADY),
  .SAXIHP1WDATA(SAXIHP1WDATA),
  .SAXIHP1WID(SAXIHP1WID),
  .SAXIHP1WLAST(SAXIHP1WLAST),
  .SAXIHP1WRISSUECAP1EN(SAXIHP1WRISSUECAP1EN),
  .SAXIHP1WSTRB(SAXIHP1WSTRB),
  .SAXIHP1WVALID(SAXIHP1WVALID),
  .SAXIHP2ACLK(SAXIHP2ACLK),
  .SAXIHP2ARADDR(SAXIHP2ARADDR),
  .SAXIHP2ARBURST(SAXIHP2ARBURST),
  .SAXIHP2ARCACHE(SAXIHP2ARCACHE),
  .SAXIHP2ARID(SAXIHP2ARID),
  .SAXIHP2ARLEN(SAXIHP2ARLEN),
  .SAXIHP2ARLOCK(SAXIHP2ARLOCK),
  .SAXIHP2ARPROT(SAXIHP2ARPROT),
  .SAXIHP2ARQOS(SAXIHP2ARQOS),
  .SAXIHP2ARSIZE(SAXIHP2ARSIZE),
  .SAXIHP2ARVALID(SAXIHP2ARVALID),
  .SAXIHP2AWADDR(SAXIHP2AWADDR),
  .SAXIHP2AWBURST(SAXIHP2AWBURST),
  .SAXIHP2AWCACHE(SAXIHP2AWCACHE),
  .SAXIHP2AWID(SAXIHP2AWID),
  .SAXIHP2AWLEN(SAXIHP2AWLEN),
  .SAXIHP2AWLOCK(SAXIHP2AWLOCK),
  .SAXIHP2AWPROT(SAXIHP2AWPROT),
  .SAXIHP2AWQOS(SAXIHP2AWQOS),
  .SAXIHP2AWSIZE(SAXIHP2AWSIZE),
  .SAXIHP2AWVALID(SAXIHP2AWVALID),
  .SAXIHP2BREADY(SAXIHP2BREADY),
  .SAXIHP2RDISSUECAP1EN(SAXIHP2RDISSUECAP1EN),
  .SAXIHP2RREADY(SAXIHP2RREADY),
  .SAXIHP2WDATA(SAXIHP2WDATA),
  .SAXIHP2WID(SAXIHP2WID),
  .SAXIHP2WLAST(SAXIHP2WLAST),
  .SAXIHP2WRISSUECAP1EN(SAXIHP2WRISSUECAP1EN),
  .SAXIHP2WSTRB(SAXIHP2WSTRB),
  .SAXIHP2WVALID(SAXIHP2WVALID),
  .SAXIHP3ACLK(SAXIHP3ACLK),
  .SAXIHP3ARADDR(SAXIHP3ARADDR),
  .SAXIHP3ARBURST(SAXIHP3ARBURST),
  .SAXIHP3ARCACHE(SAXIHP3ARCACHE),
  .SAXIHP3ARID(SAXIHP3ARID),
  .SAXIHP3ARLEN(SAXIHP3ARLEN),
  .SAXIHP3ARLOCK(SAXIHP3ARLOCK),
  .SAXIHP3ARPROT(SAXIHP3ARPROT),
  .SAXIHP3ARQOS(SAXIHP3ARQOS),
  .SAXIHP3ARSIZE(SAXIHP3ARSIZE),
  .SAXIHP3ARVALID(SAXIHP3ARVALID),
  .SAXIHP3AWADDR(SAXIHP3AWADDR),
  .SAXIHP3AWBURST(SAXIHP3AWBURST),
  .SAXIHP3AWCACHE(SAXIHP3AWCACHE),
  .SAXIHP3AWID(SAXIHP3AWID),
  .SAXIHP3AWLEN(SAXIHP3AWLEN),
  .SAXIHP3AWLOCK(SAXIHP3AWLOCK),
  .SAXIHP3AWPROT(SAXIHP3AWPROT),
  .SAXIHP3AWQOS(SAXIHP3AWQOS),
  .SAXIHP3AWSIZE(SAXIHP3AWSIZE),
  .SAXIHP3AWVALID(SAXIHP3AWVALID),
  .SAXIHP3BREADY(SAXIHP3BREADY),
  .SAXIHP3RDISSUECAP1EN(SAXIHP3RDISSUECAP1EN),
  .SAXIHP3RREADY(SAXIHP3RREADY),
  .SAXIHP3WDATA(SAXIHP3WDATA),
  .SAXIHP3WID(SAXIHP3WID),
  .SAXIHP3WLAST(SAXIHP3WLAST),
  .SAXIHP3WRISSUECAP1EN(SAXIHP3WRISSUECAP1EN),
  .SAXIHP3WSTRB(SAXIHP3WSTRB),
  .SAXIHP3WVALID(SAXIHP3WVALID)
);
// }}}

endmodule
/* vim: set fdm=marker: */
