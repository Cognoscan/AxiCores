/**
# PS7 Wrapper #

Wraps the PS7 primitive using SystemVerilog Interfaces, making for a much more 
manageable netlist.
*/
module ps7_wrapper
(
    // AXI3 Bus Masters
    axi3_if.master m_axi_gp0, ///< Master GP0 - 32-bit data, 32-bit address, 12-bit ID
    axi3_if.master m_axi_gp1, ///< Master GP0 - 32-bit data, 32-bit address, 12-bit ID

    // AXI3 ACP Bus Slave
    axi3_if.slave s_axi_acp, ///< Slave ACP - 64-bit data, 32-bit address, 3-bit ID
    input [4:0] s_axi_acp_awuser, ///< Slave ACP - User pins to inform Snoop Control Unit
    input [4:0] s_axi_acp_aruser, ///< Slave ACP - User pins to inform Snoop Control Unit

    // AXI3 Bus Slaves
    axi3_if.slave s_axi_gp0, ///< Slave GP0 - 32-bit data, 32-bit address, 6-bit ID
    axi3_if.slave s_axi_gp1, ///< Slave GP1 - 32-bit data, 32-bit address, 6-bit ID
    axi3_if.slave s_axi_hp0, ///< Slave HP0 - 64-bit data, 32-bit address, 6-bit ID
    axi3_if.slave s_axi_hp1, ///< Slave HP1 - 64-bit data, 32-bit address, 6-bit ID
    axi3_if.slave s_axi_hp2, ///< Slave HP2 - 64-bit data, 32-bit address, 6-bit ID
    axi3_if.slave s_axi_hp3, ///< Slave HP3 - 64-bit data, 32-bit address, 6-bit ID

    // AXI3 Bus Slave FIFO Interfaces
    axi_hp_fifo_if.slave s_axi_hp0_fifo, ///< Slave HP0 - FIFO Control
    axi_hp_fifo_if.slave s_axi_hp1_fifo, ///< Slave HP1 - FIFO Control
    axi_hp_fifo_if.slave s_axi_hp2_fifo, ///< Slave HP2 - FIFO Control
    axi_hp_fifo_if.slave s_axi_hp3_fifo, ///< Slave HP3 - FIFO Control

    // DMA Peripheral Request Interfaces
    dma_req_if.zynq dma0, ///< DMA0 request interface
    dma_req_if.zynq dma1, ///< DMA1 request interface
    dma_req_if.zynq dma2, ///< DMA2 request interface
    dma_req_if.zynq dma3  ///< DMA3 request interface

);

// }}}
///////////////////////////////////////////////////////////////////////////
// Signal Declarations {{{
///////////////////////////////////////////////////////////////////////////

// DDR
wire [31:0] DDRDQ; //inout
wire [14:0] DDRA; //inout
wire [3:0] DDRARB; //input
wire [3:0] DDRDM; //inout
wire [3:0] DDRDQSN; //inout
wire [3:0] DDRDQSP; //inout
wire [2:0] DDRBA; //inout
wire DDRCASB; //inout
wire DDRCKE; //inout
wire DDRCKN; //inout
wire DDRCKP; //inout
wire DDRCSB; //inout
wire DDRDRSTB; //inout
wire DDRODT; //inout
wire DDRRASB; //inout
wire DDRVRN; //inout
wire DDRVRP; //inout
wire DDRWEB; //inout

// DMA0
wire [1:0] DMA0DATYPE; //output
wire [1:0] DMA0DRTYPE; //input
wire DMA0ACLK; //input
wire DMA0DAREADY; //input
wire DMA0DAVALID; //output
wire DMA0DRLAST; //input
wire DMA0DRREADY; //output
wire DMA0DRVALID; //input
wire DMA0RSTN; //output

// DMA1
wire [1:0] DMA1DATYPE; //output
wire [1:0] DMA1DRTYPE; //input
wire DMA1ACLK; //input
wire DMA1DAREADY; //input
wire DMA1DAVALID; //output
wire DMA1DRLAST; //input
wire DMA1DRREADY; //output
wire DMA1DRVALID; //input
wire DMA1RSTN; //output

// DMA2
wire [1:0] DMA2DATYPE; //output
wire [1:0] DMA2DRTYPE; //input
wire DMA2ACLK; //input
wire DMA2DAREADY; //input
wire DMA2DAVALID; //output
wire DMA2DRLAST; //input
wire DMA2DRREADY; //output
wire DMA2DRVALID; //input
wire DMA2RSTN; //output

// DMA3
wire [1:0] DMA3DATYPE; //output
wire [1:0] DMA3DRTYPE; //input
wire DMA3ACLK; //input
wire DMA3DAREADY; //input
wire DMA3DAVALID; //output
wire DMA3DRLAST; //input
wire DMA3DRREADY; //output
wire DMA3DRVALID; //input
wire DMA3RSTN; //output

// EMIOCAN0
wire EMIOCAN0PHYRX; //input
wire EMIOCAN0PHYTX; //output

// EMIOCAN1
wire EMIOCAN1PHYRX; //input
wire EMIOCAN1PHYTX; //output

// EMIOENET0
wire [7:0] EMIOENET0GMIIRXD; //input
wire [7:0] EMIOENET0GMIITXD; //output
wire EMIOENET0EXTINTIN; //input
wire EMIOENET0GMIICOL; //input
wire EMIOENET0GMIICRS; //input
wire EMIOENET0GMIIRXCLK; //input
wire EMIOENET0GMIIRXDV; //input
wire EMIOENET0GMIIRXER; //input
wire EMIOENET0GMIITXCLK; //input
wire EMIOENET0GMIITXEN; //output
wire EMIOENET0GMIITXER; //output
wire EMIOENET0MDIOI; //input
wire EMIOENET0MDIOMDC; //output
wire EMIOENET0MDIOO; //output
wire EMIOENET0MDIOTN; //output
wire EMIOENET0PTPDELAYREQRX; //output
wire EMIOENET0PTPDELAYREQTX; //output
wire EMIOENET0PTPPDELAYREQRX; //output
wire EMIOENET0PTPPDELAYREQTX; //output
wire EMIOENET0PTPPDELAYRESPRX; //output
wire EMIOENET0PTPPDELAYRESPTX; //output
wire EMIOENET0PTPSYNCFRAMERX; //output
wire EMIOENET0PTPSYNCFRAMETX; //output
wire EMIOENET0SOFRX; //output
wire EMIOENET0SOFTX; //output

// EMIOENET1
wire [7:0] EMIOENET1GMIIRXD; //input
wire [7:0] EMIOENET1GMIITXD; //output
wire EMIOENET1EXTINTIN; //input
wire EMIOENET1GMIICOL; //input
wire EMIOENET1GMIICRS; //input
wire EMIOENET1GMIIRXCLK; //input
wire EMIOENET1GMIIRXDV; //input
wire EMIOENET1GMIIRXER; //input
wire EMIOENET1GMIITXCLK; //input
wire EMIOENET1GMIITXEN; //output
wire EMIOENET1GMIITXER; //output
wire EMIOENET1MDIOI; //input
wire EMIOENET1MDIOMDC; //output
wire EMIOENET1MDIOO; //output
wire EMIOENET1MDIOTN; //output
wire EMIOENET1PTPDELAYREQRX; //output
wire EMIOENET1PTPDELAYREQTX; //output
wire EMIOENET1PTPPDELAYREQRX; //output
wire EMIOENET1PTPPDELAYREQTX; //output
wire EMIOENET1PTPPDELAYRESPRX; //output
wire EMIOENET1PTPPDELAYRESPTX; //output
wire EMIOENET1PTPSYNCFRAMERX; //output
wire EMIOENET1PTPSYNCFRAMETX; //output
wire EMIOENET1SOFRX; //output
wire EMIOENET1SOFTX; //output

// EMIOI2C0
wire EMIOI2C0SCLI; //input
wire EMIOI2C0SCLO; //output
wire EMIOI2C0SCLTN; //output
wire EMIOI2C0SDAI; //input
wire EMIOI2C0SDAO; //output
wire EMIOI2C0SDATN; //output

// EMIOI2C1
wire EMIOI2C1SCLI; //input
wire EMIOI2C1SCLO; //output
wire EMIOI2C1SCLTN; //output
wire EMIOI2C1SDAI; //input
wire EMIOI2C1SDAO; //output
wire EMIOI2C1SDATN; //output

// EMIOPJTAG
wire EMIOPJTAGTCK; //input
wire EMIOPJTAGTDI; //input
wire EMIOPJTAGTDO; //output
wire EMIOPJTAGTDTN; //output
wire EMIOPJTAGTMS; //input

// EMIOSDIO0
wire [3:0] EMIOSDIO0DATAI; //input
wire [3:0] EMIOSDIO0DATAO; //output
wire [3:0] EMIOSDIO0DATATN; //output
wire [2:0] EMIOSDIO0BUSVOLT; //output
wire EMIOSDIO0BUSPOW; //output
wire EMIOSDIO0CDN; //input
wire EMIOSDIO0CLK; //output
wire EMIOSDIO0CLKFB; //input
wire EMIOSDIO0CMDI; //input
wire EMIOSDIO0CMDO; //output
wire EMIOSDIO0CMDTN; //output
wire EMIOSDIO0LED; //output
wire EMIOSDIO0WP; //input

// EMIOSDIO1
wire [3:0] EMIOSDIO1DATAI; //input
wire [3:0] EMIOSDIO1DATAO; //output
wire [3:0] EMIOSDIO1DATATN; //output
wire [2:0] EMIOSDIO1BUSVOLT; //output
wire EMIOSDIO1BUSPOW; //output
wire EMIOSDIO1CDN; //input
wire EMIOSDIO1CLK; //output
wire EMIOSDIO1CLKFB; //input
wire EMIOSDIO1CMDI; //input
wire EMIOSDIO1CMDO; //output
wire EMIOSDIO1CMDTN; //output
wire EMIOSDIO1LED; //output
wire EMIOSDIO1WP; //input

// EMIOSPI0
wire [2:0] EMIOSPI0SSON; //output
wire EMIOSPI0MI; //input
wire EMIOSPI0MO; //output
wire EMIOSPI0MOTN; //output
wire EMIOSPI0SCLKI; //input
wire EMIOSPI0SCLKO; //output
wire EMIOSPI0SCLKTN; //output
wire EMIOSPI0SI; //input
wire EMIOSPI0SO; //output
wire EMIOSPI0SSIN; //input
wire EMIOSPI0SSNTN; //output
wire EMIOSPI0STN; //output

// EMIOSPI1
wire [2:0] EMIOSPI1SSON; //output
wire EMIOSPI1MI; //input
wire EMIOSPI1MO; //output
wire EMIOSPI1MOTN; //output
wire EMIOSPI1SCLKI; //input
wire EMIOSPI1SCLKO; //output
wire EMIOSPI1SCLKTN; //output
wire EMIOSPI1SI; //input
wire EMIOSPI1SO; //output
wire EMIOSPI1SSIN; //input
wire EMIOSPI1SSNTN; //output
wire EMIOSPI1STN; //output

// EMIO Misc
wire EMIOSRAMINTIN; //input

// EMIOTRACE
wire [31:0] EMIOTRACEDATA; //output
wire EMIOTRACECLK; //input
wire EMIOTRACECTL; //output

// EMIOUART0
wire EMIOUART0CTSN; //input
wire EMIOUART0DCDN; //input
wire EMIOUART0DSRN; //input
wire EMIOUART0DTRN; //output
wire EMIOUART0RIN; //input
wire EMIOUART0RTSN; //output
wire EMIOUART0RX; //input
wire EMIOUART0TX; //output

// EMIOUART1
wire EMIOUART1CTSN; //input
wire EMIOUART1DCDN; //input
wire EMIOUART1DSRN; //input
wire EMIOUART1DTRN; //output
wire EMIOUART1RIN; //input
wire EMIOUART1RTSN; //output
wire EMIOUART1RX; //input
wire EMIOUART1TX; //output

// EMIOUSB0
wire [1:0] EMIOUSB0PORTINDCTL; //output
wire EMIOUSB0VBUSPWRFAULT; //input
wire EMIOUSB0VBUSPWRSELECT; //output

// EMIOUSB0
wire [1:0] EMIOUSB1PORTINDCTL; //output
wire EMIOUSB1VBUSPWRFAULT; //input
wire EMIOUSB1VBUSPWRSELECT; //output

wire EMIOWDTCLKI; //input
wire EMIOWDTRSTO; //output

// EVENT
wire [1:0] EVENTSTANDBYWFE; //output
wire [1:0] EVENTSTANDBYWFI; //output
wire EVENTEVENTI; //input
wire EVENTEVENTO; //output

wire FPGAIDLEN; //input

// FTM
wire [31:0] FTMDTRACEINDATA; //input
wire [31:0] FTMTF2PDEBUG; //input
wire [31:0] FTMTP2FDEBUG; //output
wire [3:0] FTMDTRACEINATID; //input
wire [3:0] FTMTF2PTRIG; //input
wire [3:0] FTMTF2PTRIGACK; //output
wire [3:0] FTMTP2FTRIG; //output
wire [3:0] FTMTP2FTRIGACK; //input
wire FTMDTRACEINCLOCK; //input
wire FTMDTRACEINVALID; //input

// PS
wire PSCLK; //inout
wire PSPORB; //inout
wire PSSRSTB; //inout

wire [19:0] IRQF2P; //input

wire [28:0] IRQP2F; //output

// EMIOTTC0
wire [2:0] EMIOTTC0CLKI; //input
wire [2:0] EMIOTTC0WAVEO; //output

// EMIOTTC1
wire [2:0] EMIOTTC1CLKI; //input
wire [2:0] EMIOTTC1WAVEO; //output

// FCLK
wire [3:0] FCLKCLK; //output
wire [3:0] FCLKCLKTRIGN; //input
wire [3:0] FCLKRESETN; //output

wire [53:0] MIO; //inout

// EMIOGPIO
wire [63:0] EMIOGPIOI; //input
wire [63:0] EMIOGPIOO; //output
wire [63:0] EMIOGPIOTN; //output

// }}}
///////////////////////////////////////////////////////////////////////////
// Signal Bundling into Interfaces {{{
///////////////////////////////////////////////////////////////////////////

// MAXIGP0
// MAXIGP1

// }}}
///////////////////////////////////////////////////////////////////////////
// Processor Module {{{
///////////////////////////////////////////////////////////////////////////

PS7 processor (
  .DMA0DATYPE(dma0.DATYPE),
  .DMA0DAVALID(dma0.DAVALID),
  .DMA0DRREADY(dma0.DRREADY),
  .DMA0RSTN(dma0.RSTN),
  .DMA1DATYPE(dma1.DATYPE),
  .DMA1DAVALID(dma1.DAVALID),
  .DMA1DRREADY(dma1.DRREADY),
  .DMA1RSTN(dma1.RSTN),
  .DMA2DATYPE(dma2.DATYPE),
  .DMA2DAVALID(dma2.DAVALID),
  .DMA2DRREADY(dma2.DRREADY),
  .DMA2RSTN(dma2.RSTN),
  .DMA3DATYPE(dma3.DATYPE),
  .DMA3DAVALID(dma3.DAVALID),
  .DMA3DRREADY(dma3.DRREADY),
  .DMA3RSTN(dma3.RSTN),
  .EMIOCAN0PHYTX(EMIOCAN0PHYTX),
  .EMIOCAN1PHYTX(EMIOCAN1PHYTX),
  .EMIOENET0GMIITXD(EMIOENET0GMIITXD),
  .EMIOENET0GMIITXEN(EMIOENET0GMIITXEN),
  .EMIOENET0GMIITXER(EMIOENET0GMIITXER),
  .EMIOENET0MDIOMDC(EMIOENET0MDIOMDC),
  .EMIOENET0MDIOO(EMIOENET0MDIOO),
  .EMIOENET0MDIOTN(EMIOENET0MDIOTN),
  .EMIOENET0PTPDELAYREQRX(EMIOENET0PTPDELAYREQRX),
  .EMIOENET0PTPDELAYREQTX(EMIOENET0PTPDELAYREQTX),
  .EMIOENET0PTPPDELAYREQRX(EMIOENET0PTPPDELAYREQRX),
  .EMIOENET0PTPPDELAYREQTX(EMIOENET0PTPPDELAYREQTX),
  .EMIOENET0PTPPDELAYRESPRX(EMIOENET0PTPPDELAYRESPRX),
  .EMIOENET0PTPPDELAYRESPTX(EMIOENET0PTPPDELAYRESPTX),
  .EMIOENET0PTPSYNCFRAMERX(EMIOENET0PTPSYNCFRAMERX),
  .EMIOENET0PTPSYNCFRAMETX(EMIOENET0PTPSYNCFRAMETX),
  .EMIOENET0SOFRX(EMIOENET0SOFRX),
  .EMIOENET0SOFTX(EMIOENET0SOFTX),
  .EMIOENET1GMIITXD(EMIOENET1GMIITXD),
  .EMIOENET1GMIITXEN(EMIOENET1GMIITXEN),
  .EMIOENET1GMIITXER(EMIOENET1GMIITXER),
  .EMIOENET1MDIOMDC(EMIOENET1MDIOMDC),
  .EMIOENET1MDIOO(EMIOENET1MDIOO),
  .EMIOENET1MDIOTN(EMIOENET1MDIOTN),
  .EMIOENET1PTPDELAYREQRX(EMIOENET1PTPDELAYREQRX),
  .EMIOENET1PTPDELAYREQTX(EMIOENET1PTPDELAYREQTX),
  .EMIOENET1PTPPDELAYREQRX(EMIOENET1PTPPDELAYREQRX),
  .EMIOENET1PTPPDELAYREQTX(EMIOENET1PTPPDELAYREQTX),
  .EMIOENET1PTPPDELAYRESPRX(EMIOENET1PTPPDELAYRESPRX),
  .EMIOENET1PTPPDELAYRESPTX(EMIOENET1PTPPDELAYRESPTX),
  .EMIOENET1PTPSYNCFRAMERX(EMIOENET1PTPSYNCFRAMERX),
  .EMIOENET1PTPSYNCFRAMETX(EMIOENET1PTPSYNCFRAMETX),
  .EMIOENET1SOFRX(EMIOENET1SOFRX),
  .EMIOENET1SOFTX(EMIOENET1SOFTX),
  .EMIOGPIOO(EMIOGPIOO),
  .EMIOGPIOTN(EMIOGPIOTN),
  .EMIOI2C0SCLO(EMIOI2C0SCLO),
  .EMIOI2C0SCLTN(EMIOI2C0SCLTN),
  .EMIOI2C0SDAO(EMIOI2C0SDAO),
  .EMIOI2C0SDATN(EMIOI2C0SDATN),
  .EMIOI2C1SCLO(EMIOI2C1SCLO),
  .EMIOI2C1SCLTN(EMIOI2C1SCLTN),
  .EMIOI2C1SDAO(EMIOI2C1SDAO),
  .EMIOI2C1SDATN(EMIOI2C1SDATN),
  .EMIOPJTAGTDO(EMIOPJTAGTDO),
  .EMIOPJTAGTDTN(EMIOPJTAGTDTN),
  .EMIOSDIO0BUSPOW(EMIOSDIO0BUSPOW),
  .EMIOSDIO0BUSVOLT(EMIOSDIO0BUSVOLT),
  .EMIOSDIO0CLK(EMIOSDIO0CLK),
  .EMIOSDIO0CMDO(EMIOSDIO0CMDO),
  .EMIOSDIO0CMDTN(EMIOSDIO0CMDTN),
  .EMIOSDIO0DATAO(EMIOSDIO0DATAO),
  .EMIOSDIO0DATATN(EMIOSDIO0DATATN),
  .EMIOSDIO0LED(EMIOSDIO0LED),
  .EMIOSDIO1BUSPOW(EMIOSDIO1BUSPOW),
  .EMIOSDIO1BUSVOLT(EMIOSDIO1BUSVOLT),
  .EMIOSDIO1CLK(EMIOSDIO1CLK),
  .EMIOSDIO1CMDO(EMIOSDIO1CMDO),
  .EMIOSDIO1CMDTN(EMIOSDIO1CMDTN),
  .EMIOSDIO1DATAO(EMIOSDIO1DATAO),
  .EMIOSDIO1DATATN(EMIOSDIO1DATATN),
  .EMIOSDIO1LED(EMIOSDIO1LED),
  .EMIOSPI0MO(EMIOSPI0MO),
  .EMIOSPI0MOTN(EMIOSPI0MOTN),
  .EMIOSPI0SCLKO(EMIOSPI0SCLKO),
  .EMIOSPI0SCLKTN(EMIOSPI0SCLKTN),
  .EMIOSPI0SO(EMIOSPI0SO),
  .EMIOSPI0SSNTN(EMIOSPI0SSNTN),
  .EMIOSPI0SSON(EMIOSPI0SSON),
  .EMIOSPI0STN(EMIOSPI0STN),
  .EMIOSPI1MO(EMIOSPI1MO),
  .EMIOSPI1MOTN(EMIOSPI1MOTN),
  .EMIOSPI1SCLKO(EMIOSPI1SCLKO),
  .EMIOSPI1SCLKTN(EMIOSPI1SCLKTN),
  .EMIOSPI1SO(EMIOSPI1SO),
  .EMIOSPI1SSNTN(EMIOSPI1SSNTN),
  .EMIOSPI1SSON(EMIOSPI1SSON),
  .EMIOSPI1STN(EMIOSPI1STN),
  .EMIOTRACECTL(EMIOTRACECTL),
  .EMIOTRACEDATA(EMIOTRACEDATA),
  .EMIOTTC0WAVEO(EMIOTTC0WAVEO),
  .EMIOTTC1WAVEO(EMIOTTC1WAVEO),
  .EMIOUART0DTRN(EMIOUART0DTRN),
  .EMIOUART0RTSN(EMIOUART0RTSN),
  .EMIOUART0TX(EMIOUART0TX),
  .EMIOUART1DTRN(EMIOUART1DTRN),
  .EMIOUART1RTSN(EMIOUART1RTSN),
  .EMIOUART1TX(EMIOUART1TX),
  .EMIOUSB0PORTINDCTL(EMIOUSB0PORTINDCTL),
  .EMIOUSB0VBUSPWRSELECT(EMIOUSB0VBUSPWRSELECT),
  .EMIOUSB1PORTINDCTL(EMIOUSB1PORTINDCTL),
  .EMIOUSB1VBUSPWRSELECT(EMIOUSB1VBUSPWRSELECT),
  .EMIOWDTRSTO(EMIOWDTRSTO),
  .EVENTEVENTO(EVENTEVENTO),
  .EVENTSTANDBYWFE(EVENTSTANDBYWFE),
  .EVENTSTANDBYWFI(EVENTSTANDBYWFI),
  .FCLKCLK(FCLKCLK),
  .FCLKRESETN(FCLKRESETN),
  .FTMTF2PTRIGACK(FTMTF2PTRIGACK),
  .FTMTP2FDEBUG(FTMTP2FDEBUG),
  .FTMTP2FTRIG(FTMTP2FTRIG),
  .IRQP2F(IRQP2F),
  .MAXIGP0ARADDR(m_axi_gp0.ARADDR),
  .MAXIGP0ARBURST(m_axi_gp0.ARBURST),
  .MAXIGP0ARCACHE(m_axi_gp0.ARCACHE),
  .MAXIGP0ARESETN(m_axi_gp0.ARESETn),
  .MAXIGP0ARID(m_axi_gp0.ARID),
  .MAXIGP0ARLEN(m_axi_gp0.ARLEN),
  .MAXIGP0ARLOCK(m_axi_gp0.ARLOCK),
  .MAXIGP0ARPROT(m_axi_gp0.ARPROT),
  .MAXIGP0ARQOS(m_axi_gp0.ARQOS),
  .MAXIGP0ARSIZE(m_axi_gp0.ARSIZE),
  .MAXIGP0ARVALID(m_axi_gp0.ARVALID),
  .MAXIGP0AWADDR(m_axi_gp0.AWADDR),
  .MAXIGP0AWBURST(m_axi_gp0.AWBURST),
  .MAXIGP0AWCACHE(m_axi_gp0.AWCACHE),
  .MAXIGP0AWID(m_axi_gp0.AWID),
  .MAXIGP0AWLEN(m_axi_gp0.AWLEN),
  .MAXIGP0AWLOCK(m_axi_gp0.AWLOCK),
  .MAXIGP0AWPROT(m_axi_gp0.AWPROT),
  .MAXIGP0AWQOS(m_axi_gp0.AWQOS),
  .MAXIGP0AWSIZE(m_axi_gp0.AWSIZE),
  .MAXIGP0AWVALID(m_axi_gp0.AWVALID),
  .MAXIGP0BREADY(m_axi_gp0.BREADY),
  .MAXIGP0RREADY(m_axi_gp0.RREADY),
  .MAXIGP0WDATA(m_axi_gp0.WDATA),
  .MAXIGP0WID(m_axi_gp0.WID),
  .MAXIGP0WLAST(m_axi_gp0.WLAST),
  .MAXIGP0WSTRB(m_axi_gp0.WSTRB),
  .MAXIGP0WVALID(m_axi_gp0.WVALID),
  .MAXIGP1ARADDR(m_axi_gp1.ARADDR),
  .MAXIGP1ARBURST(m_axi_gp1.ARBURST),
  .MAXIGP1ARCACHE(m_axi_gp1.ARCACHE),
  .MAXIGP1ARESETN(m_axi_gp1.ARESETn),
  .MAXIGP1ARID(m_axi_gp1.ARID),
  .MAXIGP1ARLEN(m_axi_gp1.ARLEN),
  .MAXIGP1ARLOCK(m_axi_gp1.ARLOCK),
  .MAXIGP1ARPROT(m_axi_gp1.ARPROT),
  .MAXIGP1ARQOS(m_axi_gp1.ARQOS),
  .MAXIGP1ARSIZE(m_axi_gp1.ARSIZE),
  .MAXIGP1ARVALID(m_axi_gp1.ARVALID),
  .MAXIGP1AWADDR(m_axi_gp1.AWADDR),
  .MAXIGP1AWBURST(m_axi_gp1.AWBURST),
  .MAXIGP1AWCACHE(m_axi_gp1.AWCACHE),
  .MAXIGP1AWID(m_axi_gp1.AWID),
  .MAXIGP1AWLEN(m_axi_gp1.AWLEN),
  .MAXIGP1AWLOCK(m_axi_gp1.AWLOCK),
  .MAXIGP1AWPROT(m_axi_gp1.AWPROT),
  .MAXIGP1AWQOS(m_axi_gp1.AWQOS),
  .MAXIGP1AWSIZE(m_axi_gp1.AWSIZE),
  .MAXIGP1AWVALID(m_axi_gp1.AWVALID),
  .MAXIGP1BREADY(m_axi_gp1.BREADY),
  .MAXIGP1RREADY(m_axi_gp1.RREADY),
  .MAXIGP1WDATA(m_axi_gp1.WDATA),
  .MAXIGP1WID(m_axi_gp1.WID),
  .MAXIGP1WLAST(m_axi_gp1.WLAST),
  .MAXIGP1WSTRB(m_axi_gp1.WSTRB),
  .MAXIGP1WVALID(m_axi_gp1.WVALID),
  .SAXIACPARESETN(s_axi_acp.ARESETn),
  .SAXIACPARREADY(s_axi_acp.ARREADY),
  .SAXIACPAWREADY(s_axi_acp.AWREADY),
  .SAXIACPBID(s_axi_acp.BID),
  .SAXIACPBRESP(s_axi_acp.BRESP),
  .SAXIACPBVALID(s_axi_acp.BVALID),
  .SAXIACPRDATA(s_axi_acp.RDATA),
  .SAXIACPRID(s_axi_acp.RID),
  .SAXIACPRLAST(s_axi_acp.RLAST),
  .SAXIACPRRESP(s_axi_acp.RRESP),
  .SAXIACPRVALID(s_axi_acp.RVALID),
  .SAXIACPWREADY(s_axi_acp.WREADY),
  .SAXIGP0ARESETN(s_axi_gp0.ARESETn),
  .SAXIGP0ARREADY(s_axi_gp0.ARREADY),
  .SAXIGP0AWREADY(s_axi_gp0.AWREADY),
  .SAXIGP0BID(s_axi_gp0.BID),
  .SAXIGP0BRESP(s_axi_gp0.BRESP),
  .SAXIGP0BVALID(s_axi_gp0.BVALID),
  .SAXIGP0RDATA(s_axi_gp0.RDATA),
  .SAXIGP0RID(s_axi_gp0.RID),
  .SAXIGP0RLAST(s_axi_gp0.RLAST),
  .SAXIGP0RRESP(s_axi_gp0.RRESP),
  .SAXIGP0RVALID(s_axi_gp0.RVALID),
  .SAXIGP0WREADY(s_axi_gp0.WREADY),
  .SAXIGP1ARESETN(s_axi_gp1.ARESETn),
  .SAXIGP1ARREADY(s_axi_gp1.ARREADY),
  .SAXIGP1AWREADY(s_axi_gp1.AWREADY),
  .SAXIGP1BID(s_axi_gp1.BID),
  .SAXIGP1BRESP(s_axi_gp1.BRESP),
  .SAXIGP1BVALID(s_axi_gp1.BVALID),
  .SAXIGP1RDATA(s_axi_gp1.RDATA),
  .SAXIGP1RID(s_axi_gp1.RID),
  .SAXIGP1RLAST(s_axi_gp1.RLAST),
  .SAXIGP1RRESP(s_axi_gp1.RRESP),
  .SAXIGP1RVALID(s_axi_gp1.RVALID),
  .SAXIGP1WREADY(s_axi_gp1.WREADY),
  .SAXIHP0ARESETN(s_axi_hp0.ARESETn),
  .SAXIHP0ARREADY(s_axi_hp0.ARREADY),
  .SAXIHP0AWREADY(s_axi_hp0.AWREADY),
  .SAXIHP0BID(s_axi_hp0.BID),
  .SAXIHP0BRESP(s_axi_hp0.BRESP),
  .SAXIHP0BVALID(s_axi_hp0.BVALID),
  .SAXIHP0RACOUNT(s_axi_hp0_fifo.RACOUNT),
  .SAXIHP0RCOUNT(s_axi_hp0_fifo.RCOUNT),
  .SAXIHP0RDATA(s_axi_hp0.RDATA),
  .SAXIHP0RID(s_axi_hp0.RID),
  .SAXIHP0RLAST(s_axi_hp0.RLAST),
  .SAXIHP0RRESP(s_axi_hp0.RRESP),
  .SAXIHP0RVALID(s_axi_hp0.RVALID),
  .SAXIHP0WACOUNT(s_axi_hp0_fifo.WACOUNT),
  .SAXIHP0WCOUNT(s_axi_hp0_fifo.WCOUNT),
  .SAXIHP0WREADY(s_axi_hp0.WREADY),
  .SAXIHP1ARESETN(s_axi_hp1.ARESETn),
  .SAXIHP1ARREADY(s_axi_hp1.ARREADY),
  .SAXIHP1AWREADY(s_axi_hp1.AWREADY),
  .SAXIHP1BID(s_axi_hp1.BID),
  .SAXIHP1BRESP(s_axi_hp1.BRESP),
  .SAXIHP1BVALID(s_axi_hp1.BVALID),
  .SAXIHP1RACOUNT(s_axi_hp1_fifo.RACOUNT),
  .SAXIHP1RCOUNT(s_axi_hp1_fifo.RCOUNT),
  .SAXIHP1RDATA(s_axi_hp1.RDATA),
  .SAXIHP1RID(s_axi_hp1.RID),
  .SAXIHP1RLAST(s_axi_hp1.RLAST),
  .SAXIHP1RRESP(s_axi_hp1.RRESP),
  .SAXIHP1RVALID(s_axi_hp1.RVALID),
  .SAXIHP1WACOUNT(s_axi_hp1_fifo.WACOUNT),
  .SAXIHP1WCOUNT(s_axi_hp1_fifo.WCOUNT),
  .SAXIHP1WREADY(s_axi_hp1.WREADY),
  .SAXIHP2ARESETN(s_axi_hp2.ARESETn),
  .SAXIHP2ARREADY(s_axi_hp2.ARREADY),
  .SAXIHP2AWREADY(s_axi_hp2.AWREADY),
  .SAXIHP2BID(s_axi_hp2.BID),
  .SAXIHP2BRESP(s_axi_hp2.BRESP),
  .SAXIHP2BVALID(s_axi_hp2.BVALID),
  .SAXIHP2RACOUNT(s_axi_hp2_fifo.RACOUNT),
  .SAXIHP2RCOUNT(s_axi_hp2_fifo.RCOUNT),
  .SAXIHP2RDATA(s_axi_hp2.RDATA),
  .SAXIHP2RID(s_axi_hp2.RID),
  .SAXIHP2RLAST(s_axi_hp2.RLAST),
  .SAXIHP2RRESP(s_axi_hp2.RRESP),
  .SAXIHP2RVALID(s_axi_hp2.RVALID),
  .SAXIHP2WACOUNT(s_axi_hp2_fifo.WACOUNT),
  .SAXIHP2WCOUNT(s_axi_hp2_fifo.WCOUNT),
  .SAXIHP2WREADY(s_axi_hp2.WREADY),
  .SAXIHP3ARESETN(s_axi_hp3.ARESETn),
  .SAXIHP3ARREADY(s_axi_hp3.ARREADY),
  .SAXIHP3AWREADY(s_axi_hp3.AWREADY),
  .SAXIHP3BID(s_axi_hp3.BID),
  .SAXIHP3BRESP(s_axi_hp3.BRESP),
  .SAXIHP3BVALID(s_axi_hp3.BVALID),
  .SAXIHP3RACOUNT(s_axi_hp3_fifo.RACOUNT),
  .SAXIHP3RCOUNT(s_axi_hp3_fifo.RCOUNT),
  .SAXIHP3RDATA(s_axi_hp3.RDATA),
  .SAXIHP3RID(s_axi_hp3.RID),
  .SAXIHP3RLAST(s_axi_hp3.RLAST),
  .SAXIHP3RRESP(s_axi_hp3.RRESP),
  .SAXIHP3RVALID(s_axi_hp3.RVALID),
  .SAXIHP3WACOUNT(s_axi_hp3_fifo.WACOUNT),
  .SAXIHP3WCOUNT(s_axi_hp3_fifo.WCOUNT),
  .SAXIHP3WREADY(s_axi_hp3.WREADY),

  .DDRA(DDRA),
  .DDRBA(DDRBA),
  .DDRCASB(DDRCASB),
  .DDRCKE(DDRCKE),
  .DDRCKN(DDRCKN),
  .DDRCKP(DDRCKP),
  .DDRCSB(DDRCSB),
  .DDRDM(DDRDM),
  .DDRDQ(DDRDQ),
  .DDRDQSN(DDRDQSN),
  .DDRDQSP(DDRDQSP),
  .DDRDRSTB(DDRDRSTB),
  .DDRODT(DDRODT),
  .DDRRASB(DDRRASB),
  .DDRVRN(DDRVRN),
  .DDRVRP(DDRVRP),
  .DDRWEB(DDRWEB),
  .MIO(MIO),
  .PSCLK(PSCLK),
  .PSPORB(PSPORB),
  .PSSRSTB(PSSRSTB),

  .DDRARB(DDRARB),
  .DMA0ACLK(dma0.ACLK),
  .DMA0DAREADY(dma0.DAREADY),
  .DMA0DRLAST(dma0.DRLAST),
  .DMA0DRTYPE(dma0.DRTYPE),
  .DMA0DRVALID(dma0.DRVALID),
  .DMA1ACLK(dma1.ACLK),
  .DMA1DAREADY(dma1.DAREADY),
  .DMA1DRLAST(dma1.DRLAST),
  .DMA1DRTYPE(dma1.DRTYPE),
  .DMA1DRVALID(dma1.DRVALID),
  .DMA2ACLK(dma2.ACLK),
  .DMA2DAREADY(dma2.DAREADY),
  .DMA2DRLAST(dma2.DRLAST),
  .DMA2DRTYPE(dma2.DRTYPE),
  .DMA2DRVALID(dma2.DRVALID),
  .DMA3ACLK(dma3.ACLK),
  .DMA3DAREADY(dma3.DAREADY),
  .DMA3DRLAST(dma3.DRLAST),
  .DMA3DRTYPE(dma3.DRTYPE),
  .DMA3DRVALID(dma3.DRVALID),
  .EMIOCAN0PHYRX(EMIOCAN0PHYRX),
  .EMIOCAN1PHYRX(EMIOCAN1PHYRX),
  .EMIOENET0EXTINTIN(EMIOENET0EXTINTIN),
  .EMIOENET0GMIICOL(EMIOENET0GMIICOL),
  .EMIOENET0GMIICRS(EMIOENET0GMIICRS),
  .EMIOENET0GMIIRXCLK(EMIOENET0GMIIRXCLK),
  .EMIOENET0GMIIRXD(EMIOENET0GMIIRXD),
  .EMIOENET0GMIIRXDV(EMIOENET0GMIIRXDV),
  .EMIOENET0GMIIRXER(EMIOENET0GMIIRXER),
  .EMIOENET0GMIITXCLK(EMIOENET0GMIITXCLK),
  .EMIOENET0MDIOI(EMIOENET0MDIOI),
  .EMIOENET1EXTINTIN(EMIOENET1EXTINTIN),
  .EMIOENET1GMIICOL(EMIOENET1GMIICOL),
  .EMIOENET1GMIICRS(EMIOENET1GMIICRS),
  .EMIOENET1GMIIRXCLK(EMIOENET1GMIIRXCLK),
  .EMIOENET1GMIIRXD(EMIOENET1GMIIRXD),
  .EMIOENET1GMIIRXDV(EMIOENET1GMIIRXDV),
  .EMIOENET1GMIIRXER(EMIOENET1GMIIRXER),
  .EMIOENET1GMIITXCLK(EMIOENET1GMIITXCLK),
  .EMIOENET1MDIOI(EMIOENET1MDIOI),
  .EMIOGPIOI(EMIOGPIOI),
  .EMIOI2C0SCLI(EMIOI2C0SCLI),
  .EMIOI2C0SDAI(EMIOI2C0SDAI),
  .EMIOI2C1SCLI(EMIOI2C1SCLI),
  .EMIOI2C1SDAI(EMIOI2C1SDAI),
  .EMIOPJTAGTCK(EMIOPJTAGTCK),
  .EMIOPJTAGTDI(EMIOPJTAGTDI),
  .EMIOPJTAGTMS(EMIOPJTAGTMS),
  .EMIOSDIO0CDN(EMIOSDIO0CDN),
  .EMIOSDIO0CLKFB(EMIOSDIO0CLKFB),
  .EMIOSDIO0CMDI(EMIOSDIO0CMDI),
  .EMIOSDIO0DATAI(EMIOSDIO0DATAI),
  .EMIOSDIO0WP(EMIOSDIO0WP),
  .EMIOSDIO1CDN(EMIOSDIO1CDN),
  .EMIOSDIO1CLKFB(EMIOSDIO1CLKFB),
  .EMIOSDIO1CMDI(EMIOSDIO1CMDI),
  .EMIOSDIO1DATAI(EMIOSDIO1DATAI),
  .EMIOSDIO1WP(EMIOSDIO1WP),
  .EMIOSPI0MI(EMIOSPI0MI),
  .EMIOSPI0SCLKI(EMIOSPI0SCLKI),
  .EMIOSPI0SI(EMIOSPI0SI),
  .EMIOSPI0SSIN(EMIOSPI0SSIN),
  .EMIOSPI1MI(EMIOSPI1MI),
  .EMIOSPI1SCLKI(EMIOSPI1SCLKI),
  .EMIOSPI1SI(EMIOSPI1SI),
  .EMIOSPI1SSIN(EMIOSPI1SSIN),
  .EMIOSRAMINTIN(EMIOSRAMINTIN),
  .EMIOTRACECLK(EMIOTRACECLK),
  .EMIOTTC0CLKI(EMIOTTC0CLKI),
  .EMIOTTC1CLKI(EMIOTTC1CLKI),
  .EMIOUART0CTSN(EMIOUART0CTSN),
  .EMIOUART0DCDN(EMIOUART0DCDN),
  .EMIOUART0DSRN(EMIOUART0DSRN),
  .EMIOUART0RIN(EMIOUART0RIN),
  .EMIOUART0RX(EMIOUART0RX),
  .EMIOUART1CTSN(EMIOUART1CTSN),
  .EMIOUART1DCDN(EMIOUART1DCDN),
  .EMIOUART1DSRN(EMIOUART1DSRN),
  .EMIOUART1RIN(EMIOUART1RIN),
  .EMIOUART1RX(EMIOUART1RX),
  .EMIOUSB0VBUSPWRFAULT(EMIOUSB0VBUSPWRFAULT),
  .EMIOUSB1VBUSPWRFAULT(EMIOUSB1VBUSPWRFAULT),
  .EMIOWDTCLKI(EMIOWDTCLKI),
  .EVENTEVENTI(EVENTEVENTI),
  .FCLKCLKTRIGN(FCLKCLKTRIGN),
  .FPGAIDLEN(FPGAIDLEN),
  .FTMDTRACEINATID(FTMDTRACEINATID),
  .FTMDTRACEINCLOCK(FTMDTRACEINCLOCK),
  .FTMDTRACEINDATA(FTMDTRACEINDATA),
  .FTMDTRACEINVALID(FTMDTRACEINVALID),
  .FTMTF2PDEBUG(FTMTF2PDEBUG),
  .FTMTF2PTRIG(FTMTF2PTRIG),
  .FTMTP2FTRIGACK(FTMTP2FTRIGACK),
  .IRQF2P(IRQF2P),
  .MAXIGP0ACLK(m_axi_gp0.ACLK),
  .MAXIGP0ARREADY(m_axi_gp0.ARREADY),
  .MAXIGP0AWREADY(m_axi_gp0.AWREADY),
  .MAXIGP0BID(m_axi_gp0.BID),
  .MAXIGP0BRESP(m_axi_gp0.BRESP),
  .MAXIGP0BVALID(m_axi_gp0.BVALID),
  .MAXIGP0RDATA(m_axi_gp0.RDATA),
  .MAXIGP0RID(m_axi_gp0.RID),
  .MAXIGP0RLAST(m_axi_gp0.RLAST),
  .MAXIGP0RRESP(m_axi_gp0.RRESP),
  .MAXIGP0RVALID(m_axi_gp0.RVALID),
  .MAXIGP0WREADY(m_axi_gp0.WREADY),
  .MAXIGP1ACLK(m_axi_gp1.ACLK),
  .MAXIGP1ARREADY(m_axi_gp1.ARREADY),
  .MAXIGP1AWREADY(m_axi_gp1.AWREADY),
  .MAXIGP1BID(m_axi_gp1.BID),
  .MAXIGP1BRESP(m_axi_gp1.BRESP),
  .MAXIGP1BVALID(m_axi_gp1.BVALID),
  .MAXIGP1RDATA(m_axi_gp1.RDATA),
  .MAXIGP1RID(m_axi_gp1.RID),
  .MAXIGP1RLAST(m_axi_gp1.RLAST),
  .MAXIGP1RRESP(m_axi_gp1.RRESP),
  .MAXIGP1RVALID(m_axi_gp1.RVALID),
  .MAXIGP1WREADY(m_axi_gp1.WREADY),
  .SAXIACPACLK(s_axi_acp.ACLK),
  .SAXIACPARADDR(s_axi_acp.ARADDR),
  .SAXIACPARBURST(s_axi_acp.ARBURST),
  .SAXIACPARCACHE(s_axi_acp.ARCACHE),
  .SAXIACPARID(s_axi_acp.ARID),
  .SAXIACPARLEN(s_axi_acp.ARLEN),
  .SAXIACPARLOCK(s_axi_acp.ARLOCK),
  .SAXIACPARPROT(s_axi_acp.ARPROT),
  .SAXIACPARQOS(s_axi_acp.ARQOS),
  .SAXIACPARSIZE(s_axi_acp.ARSIZE),
  .SAXIACPARUSER(s_axi_acp_aruser),
  .SAXIACPARVALID(s_axi_acp.ARVALID),
  .SAXIACPAWADDR(s_axi_acp.AWADDR),
  .SAXIACPAWBURST(s_axi_acp.AWBURST),
  .SAXIACPAWCACHE(s_axi_acp.AWCACHE),
  .SAXIACPAWID(s_axi_acp.AWID),
  .SAXIACPAWLEN(s_axi_acp.AWLEN),
  .SAXIACPAWLOCK(s_axi_acp.AWLOCK),
  .SAXIACPAWPROT(s_axi_acp.AWPROT),
  .SAXIACPAWQOS(s_axi_acp.AWQOS),
  .SAXIACPAWSIZE(s_axi_acp.AWSIZE),
  .SAXIACPAWUSER(s_axi_acp_awuser),
  .SAXIACPAWVALID(s_axi_acp.AWVALID),
  .SAXIACPBREADY(s_axi_acp.BREADY),
  .SAXIACPRREADY(s_axi_acp.RREADY),
  .SAXIACPWDATA(s_axi_acp.WDATA),
  .SAXIACPWID(s_axi_acp.WID),
  .SAXIACPWLAST(s_axi_acp.WLAST),
  .SAXIACPWSTRB(s_axi_acp.WSTRB),
  .SAXIACPWVALID(s_axi_acp.WVALID),
  .SAXIGP0ACLK(s_axi_gp0.ACLK),
  .SAXIGP0ARADDR(s_axi_gp0.ARADDR),
  .SAXIGP0ARBURST(s_axi_gp0.ARBURST),
  .SAXIGP0ARCACHE(s_axi_gp0.ARCACHE),
  .SAXIGP0ARID(s_axi_gp0.ARID),
  .SAXIGP0ARLEN(s_axi_gp0.ARLEN),
  .SAXIGP0ARLOCK(s_axi_gp0.ARLOCK),
  .SAXIGP0ARPROT(s_axi_gp0.ARPROT),
  .SAXIGP0ARQOS(s_axi_gp0.ARQOS),
  .SAXIGP0ARSIZE(s_axi_gp0.ARSIZE),
  .SAXIGP0ARVALID(s_axi_gp0.ARVALID),
  .SAXIGP0AWADDR(s_axi_gp0.AWADDR),
  .SAXIGP0AWBURST(s_axi_gp0.AWBURST),
  .SAXIGP0AWCACHE(s_axi_gp0.AWCACHE),
  .SAXIGP0AWID(s_axi_gp0.AWID),
  .SAXIGP0AWLEN(s_axi_gp0.AWLEN),
  .SAXIGP0AWLOCK(s_axi_gp0.AWLOCK),
  .SAXIGP0AWPROT(s_axi_gp0.AWPROT),
  .SAXIGP0AWQOS(s_axi_gp0.AWQOS),
  .SAXIGP0AWSIZE(s_axi_gp0.AWSIZE),
  .SAXIGP0AWVALID(s_axi_gp0.AWVALID),
  .SAXIGP0BREADY(s_axi_gp0.BREADY),
  .SAXIGP0RREADY(s_axi_gp0.RREADY),
  .SAXIGP0WDATA(s_axi_gp0.WDATA),
  .SAXIGP0WID(s_axi_gp0.WID),
  .SAXIGP0WLAST(s_axi_gp0.WLAST),
  .SAXIGP0WSTRB(s_axi_gp0.WSTRB),
  .SAXIGP0WVALID(s_axi_gp0.WVALID),
  .SAXIGP1ACLK(s_axi_gp1.ACLK),
  .SAXIGP1ARADDR(s_axi_gp1.ARADDR),
  .SAXIGP1ARBURST(s_axi_gp1.ARBURST),
  .SAXIGP1ARCACHE(s_axi_gp1.ARCACHE),
  .SAXIGP1ARID(s_axi_gp1.ARID),
  .SAXIGP1ARLEN(s_axi_gp1.ARLEN),
  .SAXIGP1ARLOCK(s_axi_gp1.ARLOCK),
  .SAXIGP1ARPROT(s_axi_gp1.ARPROT),
  .SAXIGP1ARQOS(s_axi_gp1.ARQOS),
  .SAXIGP1ARSIZE(s_axi_gp1.ARSIZE),
  .SAXIGP1ARVALID(s_axi_gp1.ARVALID),
  .SAXIGP1AWADDR(s_axi_gp1.AWADDR),
  .SAXIGP1AWBURST(s_axi_gp1.AWBURST),
  .SAXIGP1AWCACHE(s_axi_gp1.AWCACHE),
  .SAXIGP1AWID(s_axi_gp1.AWID),
  .SAXIGP1AWLEN(s_axi_gp1.AWLEN),
  .SAXIGP1AWLOCK(s_axi_gp1.AWLOCK),
  .SAXIGP1AWPROT(s_axi_gp1.AWPROT),
  .SAXIGP1AWQOS(s_axi_gp1.AWQOS),
  .SAXIGP1AWSIZE(s_axi_gp1.AWSIZE),
  .SAXIGP1AWVALID(s_axi_gp1.AWVALID),
  .SAXIGP1BREADY(s_axi_gp1.BREADY),
  .SAXIGP1RREADY(s_axi_gp1.RREADY),
  .SAXIGP1WDATA(s_axi_gp1.WDATA),
  .SAXIGP1WID(s_axi_gp1.WID),
  .SAXIGP1WLAST(s_axi_gp1.WLAST),
  .SAXIGP1WSTRB(s_axi_gp1.WSTRB),
  .SAXIGP1WVALID(s_axi_gp1.WVALID),
  .SAXIHP0ACLK(s_axi_hp0.ACLK),
  .SAXIHP0ARADDR(s_axi_hp0.ARADDR),
  .SAXIHP0ARBURST(s_axi_hp0.ARBURST),
  .SAXIHP0ARCACHE(s_axi_hp0.ARCACHE),
  .SAXIHP0ARID(s_axi_hp0.ARID),
  .SAXIHP0ARLEN(s_axi_hp0.ARLEN),
  .SAXIHP0ARLOCK(s_axi_hp0.ARLOCK),
  .SAXIHP0ARPROT(s_axi_hp0.ARPROT),
  .SAXIHP0ARQOS(s_axi_hp0.ARQOS),
  .SAXIHP0ARSIZE(s_axi_hp0.ARSIZE),
  .SAXIHP0ARVALID(s_axi_hp0.ARVALID),
  .SAXIHP0AWADDR(s_axi_hp0.AWADDR),
  .SAXIHP0AWBURST(s_axi_hp0.AWBURST),
  .SAXIHP0AWCACHE(s_axi_hp0.AWCACHE),
  .SAXIHP0AWID(s_axi_hp0.AWID),
  .SAXIHP0AWLEN(s_axi_hp0.AWLEN),
  .SAXIHP0AWLOCK(s_axi_hp0.AWLOCK),
  .SAXIHP0AWPROT(s_axi_hp0.AWPROT),
  .SAXIHP0AWQOS(s_axi_hp0.AWQOS),
  .SAXIHP0AWSIZE(s_axi_hp0.AWSIZE),
  .SAXIHP0AWVALID(s_axi_hp0.AWVALID),
  .SAXIHP0BREADY(s_axi_hp0.BREADY),
  .SAXIHP0RDISSUECAP1EN(s_axi_hp0_fifo.RDISSUECAP1EN),
  .SAXIHP0RREADY(s_axi_hp0.RREADY),
  .SAXIHP0WDATA(s_axi_hp0.WDATA),
  .SAXIHP0WID(s_axi_hp0.WID),
  .SAXIHP0WLAST(s_axi_hp0.WLAST),
  .SAXIHP0WRISSUECAP1EN(s_axi_hp0_fifo.WRISSUECAP1EN),
  .SAXIHP0WSTRB(s_axi_hp0.WSTRB),
  .SAXIHP0WVALID(s_axi_hp0.WVALID),
  .SAXIHP1ACLK(s_axi_hp1.ACLK),
  .SAXIHP1ARADDR(s_axi_hp1.ARADDR),
  .SAXIHP1ARBURST(s_axi_hp1.ARBURST),
  .SAXIHP1ARCACHE(s_axi_hp1.ARCACHE),
  .SAXIHP1ARID(s_axi_hp1.ARID),
  .SAXIHP1ARLEN(s_axi_hp1.ARLEN),
  .SAXIHP1ARLOCK(s_axi_hp1.ARLOCK),
  .SAXIHP1ARPROT(s_axi_hp1.ARPROT),
  .SAXIHP1ARQOS(s_axi_hp1.ARQOS),
  .SAXIHP1ARSIZE(s_axi_hp1.ARSIZE),
  .SAXIHP1ARVALID(s_axi_hp1.ARVALID),
  .SAXIHP1AWADDR(s_axi_hp1.AWADDR),
  .SAXIHP1AWBURST(s_axi_hp1.AWBURST),
  .SAXIHP1AWCACHE(s_axi_hp1.AWCACHE),
  .SAXIHP1AWID(s_axi_hp1.AWID),
  .SAXIHP1AWLEN(s_axi_hp1.AWLEN),
  .SAXIHP1AWLOCK(s_axi_hp1.AWLOCK),
  .SAXIHP1AWPROT(s_axi_hp1.AWPROT),
  .SAXIHP1AWQOS(s_axi_hp1.AWQOS),
  .SAXIHP1AWSIZE(s_axi_hp1.AWSIZE),
  .SAXIHP1AWVALID(s_axi_hp1.AWVALID),
  .SAXIHP1BREADY(s_axi_hp1.BREADY),
  .SAXIHP1RDISSUECAP1EN(s_axi_hp1_fifo.RDISSUECAP1EN),
  .SAXIHP1RREADY(s_axi_hp1.RREADY),
  .SAXIHP1WDATA(s_axi_hp1.WDATA),
  .SAXIHP1WID(s_axi_hp1.WID),
  .SAXIHP1WLAST(s_axi_hp1.WLAST),
  .SAXIHP1WRISSUECAP1EN(s_axi_hp1_fifo.WRISSUECAP1EN),
  .SAXIHP1WSTRB(s_axi_hp1.WSTRB),
  .SAXIHP1WVALID(s_axi_hp1.WVALID),
  .SAXIHP2ACLK(s_axi_hp2.ACLK),
  .SAXIHP2ARADDR(s_axi_hp2.ARADDR),
  .SAXIHP2ARBURST(s_axi_hp2.ARBURST),
  .SAXIHP2ARCACHE(s_axi_hp2.ARCACHE),
  .SAXIHP2ARID(s_axi_hp2.ARID),
  .SAXIHP2ARLEN(s_axi_hp2.ARLEN),
  .SAXIHP2ARLOCK(s_axi_hp2.ARLOCK),
  .SAXIHP2ARPROT(s_axi_hp2.ARPROT),
  .SAXIHP2ARQOS(s_axi_hp2.ARQOS),
  .SAXIHP2ARSIZE(s_axi_hp2.ARSIZE),
  .SAXIHP2ARVALID(s_axi_hp2.ARVALID),
  .SAXIHP2AWADDR(s_axi_hp2.AWADDR),
  .SAXIHP2AWBURST(s_axi_hp2.AWBURST),
  .SAXIHP2AWCACHE(s_axi_hp2.AWCACHE),
  .SAXIHP2AWID(s_axi_hp2.AWID),
  .SAXIHP2AWLEN(s_axi_hp2.AWLEN),
  .SAXIHP2AWLOCK(s_axi_hp2.AWLOCK),
  .SAXIHP2AWPROT(s_axi_hp2.AWPROT),
  .SAXIHP2AWQOS(s_axi_hp2.AWQOS),
  .SAXIHP2AWSIZE(s_axi_hp2.AWSIZE),
  .SAXIHP2AWVALID(s_axi_hp2.AWVALID),
  .SAXIHP2BREADY(s_axi_hp2.BREADY),
  .SAXIHP2RDISSUECAP1EN(s_axi_hp2_fifo.RDISSUECAP1EN),
  .SAXIHP2RREADY(s_axi_hp2.RREADY),
  .SAXIHP2WDATA(s_axi_hp2.WDATA),
  .SAXIHP2WID(s_axi_hp2.WID),
  .SAXIHP2WLAST(s_axi_hp2.WLAST),
  .SAXIHP2WRISSUECAP1EN(s_axi_hp2_fifo.WRISSUECAP1EN),
  .SAXIHP2WSTRB(s_axi_hp2.WSTRB),
  .SAXIHP2WVALID(s_axi_hp2.WVALID),
  .SAXIHP3ACLK(s_axi_hp3.ACLK),
  .SAXIHP3ARADDR(s_axi_hp3.ARADDR),
  .SAXIHP3ARBURST(s_axi_hp3.ARBURST),
  .SAXIHP3ARCACHE(s_axi_hp3.ARCACHE),
  .SAXIHP3ARID(s_axi_hp3.ARID),
  .SAXIHP3ARLEN(s_axi_hp3.ARLEN),
  .SAXIHP3ARLOCK(s_axi_hp3.ARLOCK),
  .SAXIHP3ARPROT(s_axi_hp3.ARPROT),
  .SAXIHP3ARQOS(s_axi_hp3.ARQOS),
  .SAXIHP3ARSIZE(s_axi_hp3.ARSIZE),
  .SAXIHP3ARVALID(s_axi_hp3.ARVALID),
  .SAXIHP3AWADDR(s_axi_hp3.AWADDR),
  .SAXIHP3AWBURST(s_axi_hp3.AWBURST),
  .SAXIHP3AWCACHE(s_axi_hp3.AWCACHE),
  .SAXIHP3AWID(s_axi_hp3.AWID),
  .SAXIHP3AWLEN(s_axi_hp3.AWLEN),
  .SAXIHP3AWLOCK(s_axi_hp3.AWLOCK),
  .SAXIHP3AWPROT(s_axi_hp3.AWPROT),
  .SAXIHP3AWQOS(s_axi_hp3.AWQOS),
  .SAXIHP3AWSIZE(s_axi_hp3.AWSIZE),
  .SAXIHP3AWVALID(s_axi_hp3.AWVALID),
  .SAXIHP3BREADY(s_axi_hp3.BREADY),
  .SAXIHP3RDISSUECAP1EN(s_axi_hp3_fifo.RDISSUECAP1EN),
  .SAXIHP3RREADY(s_axi_hp3.RREADY),
  .SAXIHP3WDATA(s_axi_hp3.WDATA),
  .SAXIHP3WID(s_axi_hp3.WID),
  .SAXIHP3WLAST(s_axi_hp3.WLAST),
  .SAXIHP3WRISSUECAP1EN(s_axi_hp3_fifo.WRISSUECAP1EN),
  .SAXIHP3WSTRB(s_axi_hp3.WSTRB),
  .SAXIHP3WVALID(s_axi_hp3.WVALID)
);
// }}}

endmodule
/* vim: set fdm=marker: */
